module aoc_solver (
    write_addr,
    write_enable,
    clear,
    clock,
    write_data,
    read_addr,
    read_data
);

    input [3:0] write_addr;
    input write_enable;
    input clear;
    input clock;
    input [31:0] write_data;
    input [3:0] read_addr;
    output [31:0] read_data;

    wire [14:0] _3891;
    wire [15:0] _3892;
    wire [15:0] _3889;
    wire [15:0] _3886;
    wire [15:0] _3883;
    wire [15:0] _3880;
    wire [15:0] _3877;
    wire [15:0] _3874;
    wire [15:0] _3871;
    wire [15:0] _3868;
    wire [15:0] _3865;
    wire [15:0] _3862;
    wire [15:0] _3859;
    wire [15:0] _3856;
    wire [15:0] _3853;
    wire [15:0] _3850;
    wire [15:0] _3847;
    wire [15:0] _3844;
    wire [15:0] _3841;
    wire [15:0] _3838;
    wire [15:0] _3835;
    wire [15:0] _3832;
    wire [15:0] _3829;
    wire [15:0] _3826;
    wire [15:0] _3823;
    wire [15:0] _3820;
    wire [15:0] _3817;
    wire [15:0] _3814;
    wire [15:0] _3811;
    wire [15:0] _3808;
    wire [15:0] _3805;
    wire [15:0] _3802;
    wire [15:0] _3799;
    wire [15:0] _3796;
    wire [15:0] _3793;
    wire [15:0] _3790;
    wire [15:0] _3787;
    wire [15:0] _3784;
    wire [15:0] _3781;
    wire [15:0] _3778;
    wire [15:0] _3775;
    wire [15:0] _3772;
    wire [15:0] _3769;
    wire [15:0] _3766;
    wire [15:0] _3763;
    wire [15:0] _3760;
    wire [15:0] _3757;
    wire [15:0] _3754;
    wire [15:0] _3751;
    wire [15:0] _3748;
    wire [15:0] _3745;
    wire [15:0] _3742;
    wire [15:0] _3739;
    wire [15:0] _3736;
    wire [15:0] _3733;
    wire [15:0] _3730;
    wire [15:0] _3727;
    wire [15:0] _3724;
    wire [15:0] _3721;
    wire [15:0] _3718;
    wire [15:0] _3715;
    wire [15:0] _3712;
    wire [15:0] _3709;
    wire [15:0] _3706;
    wire [15:0] _3703;
    wire [15:0] _3700;
    wire [15:0] _3697;
    wire [15:0] _3694;
    wire [15:0] _3691;
    wire [15:0] _3688;
    wire [15:0] _3685;
    wire [15:0] _3682;
    wire [15:0] _3679;
    wire [15:0] _3676;
    wire [15:0] _3673;
    wire [15:0] _3670;
    wire [15:0] _3667;
    wire [15:0] _3664;
    wire [15:0] _3661;
    wire [15:0] _3658;
    wire [15:0] _3655;
    wire [15:0] _3652;
    wire [15:0] _3649;
    wire [15:0] _3646;
    wire [15:0] _3643;
    wire [15:0] _3640;
    wire [15:0] _3637;
    wire [15:0] _3634;
    wire [15:0] _3631;
    wire [15:0] _3628;
    wire [15:0] _3625;
    wire [15:0] _3622;
    wire [15:0] _3619;
    wire [15:0] _3616;
    wire [15:0] _3613;
    wire [15:0] _3610;
    wire [15:0] _3607;
    wire [15:0] _3604;
    wire [15:0] _3601;
    wire [15:0] _3598;
    wire [15:0] _3596;
    wire [15:0] _3599;
    wire [15:0] _3602;
    wire [15:0] _3605;
    wire [15:0] _3608;
    wire [15:0] _3611;
    wire [15:0] _3614;
    wire [15:0] _3617;
    wire [15:0] _3620;
    wire [15:0] _3623;
    wire [15:0] _3626;
    wire [15:0] _3629;
    wire [15:0] _3632;
    wire [15:0] _3635;
    wire [15:0] _3638;
    wire [15:0] _3641;
    wire [15:0] _3644;
    wire [15:0] _3647;
    wire [15:0] _3650;
    wire [15:0] _3653;
    wire [15:0] _3656;
    wire [15:0] _3659;
    wire [15:0] _3662;
    wire [15:0] _3665;
    wire [15:0] _3668;
    wire [15:0] _3671;
    wire [15:0] _3674;
    wire [15:0] _3677;
    wire [15:0] _3680;
    wire [15:0] _3683;
    wire [15:0] _3686;
    wire [15:0] _3689;
    wire [15:0] _3692;
    wire [15:0] _3695;
    wire [15:0] _3698;
    wire [15:0] _3701;
    wire [15:0] _3704;
    wire [15:0] _3707;
    wire [15:0] _3710;
    wire [15:0] _3713;
    wire [15:0] _3716;
    wire [15:0] _3719;
    wire [15:0] _3722;
    wire [15:0] _3725;
    wire [15:0] _3728;
    wire [15:0] _3731;
    wire [15:0] _3734;
    wire [15:0] _3737;
    wire [15:0] _3740;
    wire [15:0] _3743;
    wire [15:0] _3746;
    wire [15:0] _3749;
    wire [15:0] _3752;
    wire [15:0] _3755;
    wire [15:0] _3758;
    wire [15:0] _3761;
    wire [15:0] _3764;
    wire [15:0] _3767;
    wire [15:0] _3770;
    wire [15:0] _3773;
    wire [15:0] _3776;
    wire [15:0] _3779;
    wire [15:0] _3782;
    wire [15:0] _3785;
    wire [15:0] _3788;
    wire [15:0] _3791;
    wire [15:0] _3794;
    wire [15:0] _3797;
    wire [15:0] _3800;
    wire [15:0] _3803;
    wire [15:0] _3806;
    wire [15:0] _3809;
    wire [15:0] _3812;
    wire [15:0] _3815;
    wire [15:0] _3818;
    wire [15:0] _3821;
    wire [15:0] _3824;
    wire [15:0] _3827;
    wire [15:0] _3830;
    wire [15:0] _3833;
    wire [15:0] _3836;
    wire [15:0] _3839;
    wire [15:0] _3842;
    wire [15:0] _3845;
    wire [15:0] _3848;
    wire [15:0] _3851;
    wire [15:0] _3854;
    wire [15:0] _3857;
    wire [15:0] _3860;
    wire [15:0] _3863;
    wire [15:0] _3866;
    wire [15:0] _3869;
    wire [15:0] _3872;
    wire [15:0] _3875;
    wire [15:0] _3878;
    wire [15:0] _3881;
    wire [15:0] _3884;
    wire [15:0] _3887;
    wire [15:0] _3890;
    wire [15:0] _3893;
    wire [15:0] _3594;
    wire [31:0] _3894;
    wire [15:0] _527;
    wire [15:0] _227;
    wire [15:0] _528;
    wire [15:0] _1;
    reg [15:0] _225;
    wire [31:0] _3593;
    wire _552;
    wire _553;
    wire _2;
    wire [15:0] _525;
    wire _575;
    wire _576;
    wire _3;
    wire [15:0] _522;
    wire _598;
    wire _599;
    wire _4;
    wire [15:0] _519;
    wire _621;
    wire _622;
    wire _5;
    wire [15:0] _516;
    wire _644;
    wire _645;
    wire _6;
    wire [15:0] _513;
    wire _667;
    wire _668;
    wire _7;
    wire [15:0] _510;
    wire _690;
    wire _691;
    wire _8;
    wire [15:0] _507;
    wire _713;
    wire _714;
    wire _9;
    wire [15:0] _504;
    wire _736;
    wire _737;
    wire _10;
    wire [15:0] _501;
    wire _749;
    wire _750;
    wire _11;
    wire [15:0] _498;
    wire _772;
    wire _773;
    wire _12;
    wire [15:0] _495;
    wire _802;
    wire _803;
    wire _13;
    wire [15:0] _492;
    wire _832;
    wire _833;
    wire _14;
    wire [15:0] _489;
    wire _862;
    wire _863;
    wire _15;
    wire [15:0] _486;
    wire _892;
    wire _893;
    wire _16;
    wire [15:0] _483;
    wire _922;
    wire _923;
    wire _17;
    wire [15:0] _480;
    wire _952;
    wire _953;
    wire _18;
    wire [15:0] _477;
    wire _982;
    wire _983;
    wire _19;
    wire [15:0] _474;
    wire _1012;
    wire _1013;
    wire _20;
    wire [15:0] _471;
    wire _1031;
    wire _1032;
    wire _21;
    wire [15:0] _468;
    wire _1054;
    wire _1055;
    wire _22;
    wire [15:0] _465;
    wire _1084;
    wire _1085;
    wire _23;
    wire [15:0] _462;
    wire _1114;
    wire _1115;
    wire _24;
    wire [15:0] _459;
    wire _1144;
    wire _1145;
    wire _25;
    wire [15:0] _456;
    wire _1174;
    wire _1175;
    wire _26;
    wire [15:0] _453;
    wire _1204;
    wire _1205;
    wire _27;
    wire [15:0] _450;
    wire _1234;
    wire _1235;
    wire _28;
    wire [15:0] _447;
    wire _1264;
    wire _1265;
    wire _29;
    wire [15:0] _444;
    wire _1294;
    wire _1295;
    wire _30;
    wire [15:0] _441;
    wire _1313;
    wire _1314;
    wire _31;
    wire [15:0] _438;
    wire _1336;
    wire _1337;
    wire _32;
    wire [15:0] _435;
    wire _1366;
    wire _1367;
    wire _33;
    wire [15:0] _432;
    wire _1396;
    wire _1397;
    wire _34;
    wire [15:0] _429;
    wire _1426;
    wire _1427;
    wire _35;
    wire [15:0] _426;
    wire _1456;
    wire _1457;
    wire _36;
    wire [15:0] _423;
    wire _1486;
    wire _1487;
    wire _37;
    wire [15:0] _420;
    wire _1516;
    wire _1517;
    wire _38;
    wire [15:0] _417;
    wire _1546;
    wire _1547;
    wire _39;
    wire [15:0] _414;
    wire _1576;
    wire _1577;
    wire _40;
    wire [15:0] _411;
    wire _1595;
    wire _1596;
    wire _41;
    wire [15:0] _408;
    wire _1618;
    wire _1619;
    wire _42;
    wire [15:0] _405;
    wire _1648;
    wire _1649;
    wire _43;
    wire [15:0] _402;
    wire _1678;
    wire _1679;
    wire _44;
    wire [15:0] _399;
    wire _1708;
    wire _1709;
    wire _45;
    wire [15:0] _396;
    wire _1738;
    wire _1739;
    wire _46;
    wire [15:0] _393;
    wire _1768;
    wire _1769;
    wire _47;
    wire [15:0] _390;
    wire _1798;
    wire _1799;
    wire _48;
    wire [15:0] _387;
    wire _1828;
    wire _1829;
    wire _49;
    wire [15:0] _384;
    wire _1858;
    wire _1859;
    wire _50;
    wire [15:0] _381;
    wire _1877;
    wire _1878;
    wire _51;
    wire [15:0] _378;
    wire _1900;
    wire _1901;
    wire _52;
    wire [15:0] _375;
    wire _1930;
    wire _1931;
    wire _53;
    wire [15:0] _372;
    wire _1960;
    wire _1961;
    wire _54;
    wire [15:0] _369;
    wire _1990;
    wire _1991;
    wire _55;
    wire [15:0] _366;
    wire _2020;
    wire _2021;
    wire _56;
    wire [15:0] _363;
    wire _2050;
    wire _2051;
    wire _57;
    wire [15:0] _360;
    wire _2080;
    wire _2081;
    wire _58;
    wire [15:0] _357;
    wire _2110;
    wire _2111;
    wire _59;
    wire [15:0] _354;
    wire _2140;
    wire _2141;
    wire _60;
    wire [15:0] _351;
    wire _2159;
    wire _2160;
    wire _61;
    wire [15:0] _348;
    wire _2182;
    wire _2183;
    wire _62;
    wire [15:0] _345;
    wire _2212;
    wire _2213;
    wire _63;
    wire [15:0] _342;
    wire _2242;
    wire _2243;
    wire _64;
    wire [15:0] _339;
    wire _2272;
    wire _2273;
    wire _65;
    wire [15:0] _336;
    wire _2302;
    wire _2303;
    wire _66;
    wire [15:0] _333;
    wire _2332;
    wire _2333;
    wire _67;
    wire [15:0] _330;
    wire _2362;
    wire _2363;
    wire _68;
    wire [15:0] _327;
    wire _2392;
    wire _2393;
    wire _69;
    wire [15:0] _324;
    wire _2422;
    wire _2423;
    wire _70;
    wire [15:0] _321;
    wire _2441;
    wire _2442;
    wire _71;
    wire [15:0] _318;
    wire _2464;
    wire _2465;
    wire _72;
    wire [15:0] _315;
    wire _2494;
    wire _2495;
    wire _73;
    wire [15:0] _312;
    wire _2524;
    wire _2525;
    wire _74;
    wire [15:0] _309;
    wire _2554;
    wire _2555;
    wire _75;
    wire [15:0] _306;
    wire _2584;
    wire _2585;
    wire _76;
    wire [15:0] _303;
    wire _2614;
    wire _2615;
    wire _77;
    wire [15:0] _300;
    wire _2644;
    wire _2645;
    wire _78;
    wire [15:0] _297;
    wire _2674;
    wire _2675;
    wire _79;
    wire [15:0] _294;
    wire _2704;
    wire _2705;
    wire _80;
    wire [15:0] _291;
    wire _2723;
    wire _2724;
    wire _81;
    wire [15:0] _288;
    wire _2746;
    wire _2747;
    wire _82;
    wire [15:0] _285;
    wire _2776;
    wire _2777;
    wire _83;
    wire [15:0] _282;
    wire _2806;
    wire _2807;
    wire _84;
    wire [15:0] _279;
    wire _2836;
    wire _2837;
    wire _85;
    wire [15:0] _276;
    wire _2866;
    wire _2867;
    wire _86;
    wire [15:0] _273;
    wire _2896;
    wire _2897;
    wire _87;
    wire [15:0] _270;
    wire _2926;
    wire _2927;
    wire _88;
    wire [15:0] _267;
    wire _2956;
    wire _2957;
    wire _89;
    wire [15:0] _264;
    wire _2986;
    wire _2987;
    wire _90;
    wire [15:0] _261;
    wire _3005;
    wire _3006;
    wire _91;
    wire [15:0] _258;
    wire _3018;
    wire _3019;
    wire _92;
    wire [15:0] _255;
    wire _3037;
    wire _3038;
    wire _93;
    wire [15:0] _252;
    wire _3056;
    wire _3057;
    wire _94;
    wire [15:0] _249;
    wire _3075;
    wire _3076;
    wire _95;
    wire [15:0] _246;
    wire _3094;
    wire _3095;
    wire _96;
    wire [15:0] _243;
    wire _3113;
    wire _3114;
    wire _97;
    wire [15:0] _240;
    wire _3132;
    wire _3133;
    wire _98;
    wire [15:0] _237;
    wire _3151;
    wire _3152;
    wire _99;
    wire [15:0] _234;
    wire _3170;
    wire _3171;
    wire _100;
    wire [15:0] _231;
    wire [3:0] _3576;
    wire [2:0] _3573;
    wire [3:0] _3574;
    wire [3:0] _3571;
    wire _2929;
    wire [3:0] _3165;
    wire [3:0] _3162;
    wire [3:0] _3159;
    wire [3:0] _3146;
    wire [3:0] _3143;
    wire [3:0] _3140;
    wire [3:0] _3127;
    wire [3:0] _3124;
    wire [3:0] _3121;
    wire [3:0] _3108;
    wire [3:0] _3105;
    wire [3:0] _3102;
    wire [3:0] _3089;
    wire [3:0] _3086;
    wire [3:0] _3083;
    wire [3:0] _3070;
    wire [3:0] _3067;
    wire [3:0] _3064;
    wire [3:0] _3051;
    wire [3:0] _3048;
    wire [3:0] _3045;
    wire [3:0] _3032;
    wire [3:0] _3029;
    wire [3:0] _3026;
    wire [3:0] _3013;
    wire [3:0] _2771;
    wire [3:0] _2768;
    wire [3:0] _2765;
    wire [3:0] _2762;
    wire [3:0] _2801;
    wire [3:0] _2798;
    wire [3:0] _2795;
    wire [3:0] _2792;
    wire [3:0] _2831;
    wire [3:0] _2828;
    wire [3:0] _2825;
    wire [3:0] _2822;
    wire [3:0] _2861;
    wire [3:0] _2858;
    wire [3:0] _2855;
    wire [3:0] _2852;
    wire [3:0] _2891;
    wire [3:0] _2888;
    wire [3:0] _2885;
    wire [3:0] _2882;
    wire [3:0] _2921;
    wire [3:0] _2918;
    wire [3:0] _2915;
    wire [3:0] _2912;
    wire [3:0] _2951;
    wire [3:0] _2948;
    wire [3:0] _2945;
    wire [3:0] _2942;
    wire [3:0] _2981;
    wire [3:0] _2978;
    wire [3:0] _2975;
    wire [3:0] _2972;
    wire [3:0] _3000;
    wire [3:0] _2718;
    wire [3:0] _2715;
    wire [3:0] _2699;
    wire [3:0] _2696;
    wire [3:0] _2693;
    wire [3:0] _2669;
    wire [3:0] _2666;
    wire [3:0] _2663;
    wire [3:0] _2639;
    wire [3:0] _2636;
    wire [3:0] _2633;
    wire [3:0] _2609;
    wire [3:0] _2606;
    wire [3:0] _2603;
    wire [3:0] _2579;
    wire [3:0] _2576;
    wire [3:0] _2573;
    wire [3:0] _2549;
    wire [3:0] _2546;
    wire [3:0] _2543;
    wire [3:0] _2519;
    wire [3:0] _2516;
    wire [3:0] _2513;
    wire [3:0] _2489;
    wire [3:0] _2486;
    wire [3:0] _2483;
    wire [3:0] _2480;
    wire [3:0] _2477;
    wire [3:0] _2459;
    wire [3:0] _2207;
    wire [3:0] _2204;
    wire [3:0] _2201;
    wire [3:0] _2198;
    wire [3:0] _2237;
    wire [3:0] _2234;
    wire [3:0] _2231;
    wire [3:0] _2228;
    wire [3:0] _2267;
    wire [3:0] _2264;
    wire [3:0] _2261;
    wire [3:0] _2258;
    wire [3:0] _2297;
    wire [3:0] _2294;
    wire [3:0] _2291;
    wire [3:0] _2288;
    wire [3:0] _2327;
    wire [3:0] _2324;
    wire [3:0] _2321;
    wire [3:0] _2318;
    wire [3:0] _2357;
    wire [3:0] _2354;
    wire [3:0] _2351;
    wire [3:0] _2348;
    wire [3:0] _2387;
    wire [3:0] _2384;
    wire [3:0] _2381;
    wire [3:0] _2378;
    wire [3:0] _2417;
    wire [3:0] _2414;
    wire [3:0] _2411;
    wire [3:0] _2408;
    wire [3:0] _2436;
    wire [3:0] _2154;
    wire [3:0] _2151;
    wire [3:0] _2135;
    wire [3:0] _2132;
    wire [3:0] _2129;
    wire [3:0] _2105;
    wire [3:0] _2102;
    wire [3:0] _2099;
    wire [3:0] _2075;
    wire [3:0] _2072;
    wire [3:0] _2069;
    wire [3:0] _2045;
    wire [3:0] _2042;
    wire [3:0] _2039;
    wire [3:0] _2015;
    wire [3:0] _2012;
    wire [3:0] _2009;
    wire [3:0] _1985;
    wire [3:0] _1982;
    wire [3:0] _1979;
    wire [3:0] _1955;
    wire [3:0] _1952;
    wire [3:0] _1949;
    wire [3:0] _1925;
    wire [3:0] _1922;
    wire [3:0] _1919;
    wire [3:0] _1916;
    wire [3:0] _1913;
    wire [3:0] _1895;
    wire [3:0] _1643;
    wire [3:0] _1640;
    wire [3:0] _1637;
    wire [3:0] _1634;
    wire [3:0] _1673;
    wire [3:0] _1670;
    wire [3:0] _1667;
    wire [3:0] _1664;
    wire [3:0] _1703;
    wire [3:0] _1700;
    wire [3:0] _1697;
    wire [3:0] _1694;
    wire [3:0] _1733;
    wire [3:0] _1730;
    wire [3:0] _1727;
    wire [3:0] _1724;
    wire [3:0] _1763;
    wire [3:0] _1760;
    wire [3:0] _1757;
    wire [3:0] _1754;
    wire [3:0] _1793;
    wire [3:0] _1790;
    wire [3:0] _1787;
    wire [3:0] _1784;
    wire [3:0] _1823;
    wire [3:0] _1820;
    wire [3:0] _1817;
    wire [3:0] _1814;
    wire [3:0] _1853;
    wire [3:0] _1850;
    wire [3:0] _1847;
    wire [3:0] _1844;
    wire [3:0] _1872;
    wire [3:0] _1590;
    wire [3:0] _1587;
    wire [3:0] _1571;
    wire [3:0] _1568;
    wire [3:0] _1565;
    wire [3:0] _1541;
    wire [3:0] _1538;
    wire [3:0] _1535;
    wire [3:0] _1511;
    wire [3:0] _1508;
    wire [3:0] _1505;
    wire [3:0] _1481;
    wire [3:0] _1478;
    wire [3:0] _1475;
    wire [3:0] _1451;
    wire [3:0] _1448;
    wire [3:0] _1445;
    wire [3:0] _1421;
    wire [3:0] _1418;
    wire [3:0] _1415;
    wire [3:0] _1391;
    wire [3:0] _1388;
    wire [3:0] _1385;
    wire [3:0] _1361;
    wire [3:0] _1358;
    wire [3:0] _1355;
    wire [3:0] _1352;
    wire [3:0] _1349;
    wire [3:0] _1331;
    wire [3:0] _1079;
    wire [3:0] _1076;
    wire [3:0] _1073;
    wire [3:0] _1070;
    wire [3:0] _1109;
    wire [3:0] _1106;
    wire [3:0] _1103;
    wire [3:0] _1100;
    wire [3:0] _1139;
    wire [3:0] _1136;
    wire [3:0] _1133;
    wire [3:0] _1130;
    wire [3:0] _1169;
    wire [3:0] _1166;
    wire [3:0] _1163;
    wire [3:0] _1160;
    wire [3:0] _1199;
    wire [3:0] _1196;
    wire [3:0] _1193;
    wire [3:0] _1190;
    wire [3:0] _1229;
    wire [3:0] _1226;
    wire [3:0] _1223;
    wire [3:0] _1220;
    wire [3:0] _1259;
    wire [3:0] _1256;
    wire [3:0] _1253;
    wire [3:0] _1250;
    wire [3:0] _1289;
    wire [3:0] _1286;
    wire [3:0] _1283;
    wire [3:0] _1280;
    wire [3:0] _1308;
    wire [3:0] _1026;
    wire [3:0] _1023;
    wire [3:0] _1007;
    wire [3:0] _1004;
    wire [3:0] _1001;
    wire [3:0] _977;
    wire [3:0] _974;
    wire [3:0] _971;
    wire [3:0] _947;
    wire [3:0] _944;
    wire [3:0] _941;
    wire [3:0] _917;
    wire [3:0] _914;
    wire [3:0] _911;
    wire [3:0] _887;
    wire [3:0] _884;
    wire [3:0] _881;
    wire [3:0] _857;
    wire [3:0] _854;
    wire [3:0] _851;
    wire [3:0] _827;
    wire [3:0] _824;
    wire [3:0] _821;
    wire [3:0] _797;
    wire [3:0] _794;
    wire [3:0] _791;
    wire [3:0] _788;
    wire [3:0] _785;
    wire [3:0] _767;
    wire [3:0] _547;
    wire [3:0] _542;
    wire [3:0] _538;
    wire [3:0] _543;
    wire [3:0] _548;
    wire _550;
    wire _551;
    wire _3172;
    wire _3173;
    wire _3174;
    wire _3175;
    wire _101;
    reg _534;
    wire [3:0] _570;
    wire [3:0] _593;
    wire [3:0] _616;
    wire [3:0] _639;
    wire [3:0] _662;
    wire [3:0] _685;
    wire [3:0] _708;
    wire [3:0] _731;
    wire [3:0] _744;
    wire [3:0] _741;
    wire [3:0] _739;
    wire [3:0] _742;
    wire [3:0] _745;
    wire _747;
    wire _748;
    wire _3176;
    wire _3177;
    wire _3178;
    wire _3179;
    wire _102;
    reg _727;
    wire [3:0] _728;
    wire [3:0] _723;
    wire [3:0] _720;
    wire [3:0] _718;
    wire [3:0] _721;
    wire [3:0] _724;
    wire [3:0] _729;
    wire [3:0] _732;
    wire _734;
    wire _735;
    wire _3180;
    wire _3181;
    wire _3182;
    wire _3183;
    wire _103;
    reg _704;
    wire [3:0] _705;
    wire [3:0] _700;
    wire [3:0] _697;
    wire [3:0] _695;
    wire [3:0] _698;
    wire [3:0] _701;
    wire [3:0] _706;
    wire [3:0] _709;
    wire _711;
    wire _712;
    wire _3184;
    wire _3185;
    wire _3186;
    wire _3187;
    wire _104;
    reg _681;
    wire [3:0] _682;
    wire [3:0] _677;
    wire [3:0] _674;
    wire [3:0] _672;
    wire [3:0] _675;
    wire [3:0] _678;
    wire [3:0] _683;
    wire [3:0] _686;
    wire _688;
    wire _689;
    wire _3188;
    wire _3189;
    wire _3190;
    wire _3191;
    wire _105;
    reg _658;
    wire [3:0] _659;
    wire [3:0] _654;
    wire [3:0] _651;
    wire [3:0] _649;
    wire [3:0] _652;
    wire [3:0] _655;
    wire [3:0] _660;
    wire [3:0] _663;
    wire _665;
    wire _666;
    wire _3192;
    wire _3193;
    wire _3194;
    wire _3195;
    wire _106;
    reg _635;
    wire [3:0] _636;
    wire [3:0] _631;
    wire [3:0] _628;
    wire [3:0] _626;
    wire [3:0] _629;
    wire [3:0] _632;
    wire [3:0] _637;
    wire [3:0] _640;
    wire _642;
    wire _643;
    wire _3196;
    wire _3197;
    wire _3198;
    wire _3199;
    wire _107;
    reg _612;
    wire [3:0] _613;
    wire [3:0] _608;
    wire [3:0] _605;
    wire [3:0] _603;
    wire [3:0] _606;
    wire [3:0] _609;
    wire [3:0] _614;
    wire [3:0] _617;
    wire _619;
    wire _620;
    wire _3200;
    wire _3201;
    wire _3202;
    wire _3203;
    wire _108;
    reg _589;
    wire [3:0] _590;
    wire [3:0] _585;
    wire [3:0] _582;
    wire [3:0] _580;
    wire [3:0] _583;
    wire [3:0] _586;
    wire [3:0] _591;
    wire [3:0] _594;
    wire _596;
    wire _597;
    wire _3204;
    wire _3205;
    wire _3206;
    wire _3207;
    wire _109;
    reg _566;
    wire [3:0] _567;
    wire [3:0] _562;
    wire [3:0] _559;
    wire [3:0] _557;
    wire [3:0] _560;
    wire [3:0] _563;
    wire [3:0] _568;
    wire [3:0] _571;
    wire _573;
    wire _574;
    wire _3208;
    wire _3209;
    wire _3210;
    wire _3211;
    wire _110;
    reg _546;
    wire [3:0] _764;
    wire [3:0] _761;
    wire [3:0] _758;
    wire [3:0] _754;
    wire [3:0] _759;
    wire [3:0] _762;
    wire [3:0] _765;
    wire [3:0] _768;
    wire _770;
    wire _771;
    wire _3212;
    wire _3213;
    wire _3214;
    wire _3215;
    wire _111;
    reg _541;
    wire [3:0] _1049;
    wire [3:0] _1046;
    wire [3:0] _1043;
    wire [3:0] _1040;
    wire [3:0] _1036;
    wire [3:0] _1041;
    wire [3:0] _1044;
    wire [3:0] _1047;
    wire [3:0] _1050;
    wire _1052;
    wire _1053;
    wire _3216;
    wire _3217;
    wire _3218;
    wire _3219;
    wire _112;
    reg _757;
    wire [3:0] _782;
    wire [3:0] _779;
    wire [3:0] _777;
    wire [3:0] _780;
    wire [3:0] _783;
    wire [3:0] _786;
    wire [3:0] _789;
    wire [3:0] _792;
    wire [3:0] _795;
    wire [3:0] _798;
    wire _800;
    wire _801;
    wire _3220;
    wire _3221;
    wire _3222;
    wire _3223;
    wire _113;
    reg _537;
    wire [3:0] _818;
    wire [3:0] _815;
    wire [3:0] _812;
    wire [3:0] _809;
    wire [3:0] _807;
    wire [3:0] _810;
    wire [3:0] _813;
    wire [3:0] _816;
    wire [3:0] _819;
    wire [3:0] _822;
    wire [3:0] _825;
    wire [3:0] _828;
    wire _830;
    wire _831;
    wire _3224;
    wire _3225;
    wire _3226;
    wire _3227;
    wire _114;
    reg _556;
    wire [3:0] _848;
    wire [3:0] _845;
    wire [3:0] _842;
    wire [3:0] _839;
    wire [3:0] _837;
    wire [3:0] _840;
    wire [3:0] _843;
    wire [3:0] _846;
    wire [3:0] _849;
    wire [3:0] _852;
    wire [3:0] _855;
    wire [3:0] _858;
    wire _860;
    wire _861;
    wire _3228;
    wire _3229;
    wire _3230;
    wire _3231;
    wire _115;
    reg _579;
    wire [3:0] _878;
    wire [3:0] _875;
    wire [3:0] _872;
    wire [3:0] _869;
    wire [3:0] _867;
    wire [3:0] _870;
    wire [3:0] _873;
    wire [3:0] _876;
    wire [3:0] _879;
    wire [3:0] _882;
    wire [3:0] _885;
    wire [3:0] _888;
    wire _890;
    wire _891;
    wire _3232;
    wire _3233;
    wire _3234;
    wire _3235;
    wire _116;
    reg _602;
    wire [3:0] _908;
    wire [3:0] _905;
    wire [3:0] _902;
    wire [3:0] _899;
    wire [3:0] _897;
    wire [3:0] _900;
    wire [3:0] _903;
    wire [3:0] _906;
    wire [3:0] _909;
    wire [3:0] _912;
    wire [3:0] _915;
    wire [3:0] _918;
    wire _920;
    wire _921;
    wire _3236;
    wire _3237;
    wire _3238;
    wire _3239;
    wire _117;
    reg _625;
    wire [3:0] _938;
    wire [3:0] _935;
    wire [3:0] _932;
    wire [3:0] _929;
    wire [3:0] _927;
    wire [3:0] _930;
    wire [3:0] _933;
    wire [3:0] _936;
    wire [3:0] _939;
    wire [3:0] _942;
    wire [3:0] _945;
    wire [3:0] _948;
    wire _950;
    wire _951;
    wire _3240;
    wire _3241;
    wire _3242;
    wire _3243;
    wire _118;
    reg _648;
    wire [3:0] _968;
    wire [3:0] _965;
    wire [3:0] _962;
    wire [3:0] _959;
    wire [3:0] _957;
    wire [3:0] _960;
    wire [3:0] _963;
    wire [3:0] _966;
    wire [3:0] _969;
    wire [3:0] _972;
    wire [3:0] _975;
    wire [3:0] _978;
    wire _980;
    wire _981;
    wire _3244;
    wire _3245;
    wire _3246;
    wire _3247;
    wire _119;
    reg _671;
    wire [3:0] _998;
    wire [3:0] _995;
    wire [3:0] _992;
    wire [3:0] _989;
    wire [3:0] _987;
    wire [3:0] _990;
    wire [3:0] _993;
    wire [3:0] _996;
    wire [3:0] _999;
    wire [3:0] _1002;
    wire [3:0] _1005;
    wire [3:0] _1008;
    wire _1010;
    wire _1011;
    wire _3248;
    wire _3249;
    wire _3250;
    wire _3251;
    wire _120;
    reg _694;
    wire [3:0] _1020;
    wire [3:0] _1017;
    wire [3:0] _1015;
    wire [3:0] _1018;
    wire [3:0] _1021;
    wire [3:0] _1024;
    wire [3:0] _1027;
    wire _1029;
    wire _1030;
    wire _3252;
    wire _3253;
    wire _3254;
    wire _3255;
    wire _121;
    reg _717;
    wire [3:0] _1305;
    wire [3:0] _1302;
    wire [3:0] _1299;
    wire [3:0] _1297;
    wire [3:0] _1300;
    wire [3:0] _1303;
    wire [3:0] _1306;
    wire [3:0] _1309;
    wire _1311;
    wire _1312;
    wire _3256;
    wire _3257;
    wire _3258;
    wire _3259;
    wire _122;
    reg _986;
    wire [3:0] _1277;
    wire [3:0] _1274;
    wire [3:0] _1271;
    wire [3:0] _1269;
    wire [3:0] _1272;
    wire [3:0] _1275;
    wire [3:0] _1278;
    wire [3:0] _1281;
    wire [3:0] _1284;
    wire [3:0] _1287;
    wire [3:0] _1290;
    wire _1292;
    wire _1293;
    wire _3260;
    wire _3261;
    wire _3262;
    wire _3263;
    wire _123;
    reg _956;
    wire [3:0] _1247;
    wire [3:0] _1244;
    wire [3:0] _1241;
    wire [3:0] _1239;
    wire [3:0] _1242;
    wire [3:0] _1245;
    wire [3:0] _1248;
    wire [3:0] _1251;
    wire [3:0] _1254;
    wire [3:0] _1257;
    wire [3:0] _1260;
    wire _1262;
    wire _1263;
    wire _3264;
    wire _3265;
    wire _3266;
    wire _3267;
    wire _124;
    reg _926;
    wire [3:0] _1217;
    wire [3:0] _1214;
    wire [3:0] _1211;
    wire [3:0] _1209;
    wire [3:0] _1212;
    wire [3:0] _1215;
    wire [3:0] _1218;
    wire [3:0] _1221;
    wire [3:0] _1224;
    wire [3:0] _1227;
    wire [3:0] _1230;
    wire _1232;
    wire _1233;
    wire _3268;
    wire _3269;
    wire _3270;
    wire _3271;
    wire _125;
    reg _896;
    wire [3:0] _1187;
    wire [3:0] _1184;
    wire [3:0] _1181;
    wire [3:0] _1179;
    wire [3:0] _1182;
    wire [3:0] _1185;
    wire [3:0] _1188;
    wire [3:0] _1191;
    wire [3:0] _1194;
    wire [3:0] _1197;
    wire [3:0] _1200;
    wire _1202;
    wire _1203;
    wire _3272;
    wire _3273;
    wire _3274;
    wire _3275;
    wire _126;
    reg _866;
    wire [3:0] _1157;
    wire [3:0] _1154;
    wire [3:0] _1151;
    wire [3:0] _1149;
    wire [3:0] _1152;
    wire [3:0] _1155;
    wire [3:0] _1158;
    wire [3:0] _1161;
    wire [3:0] _1164;
    wire [3:0] _1167;
    wire [3:0] _1170;
    wire _1172;
    wire _1173;
    wire _3276;
    wire _3277;
    wire _3278;
    wire _3279;
    wire _127;
    reg _836;
    wire [3:0] _1127;
    wire [3:0] _1124;
    wire [3:0] _1121;
    wire [3:0] _1119;
    wire [3:0] _1122;
    wire [3:0] _1125;
    wire [3:0] _1128;
    wire [3:0] _1131;
    wire [3:0] _1134;
    wire [3:0] _1137;
    wire [3:0] _1140;
    wire _1142;
    wire _1143;
    wire _3280;
    wire _3281;
    wire _3282;
    wire _3283;
    wire _128;
    reg _806;
    wire [3:0] _1097;
    wire [3:0] _1094;
    wire [3:0] _1091;
    wire [3:0] _1089;
    wire [3:0] _1092;
    wire [3:0] _1095;
    wire [3:0] _1098;
    wire [3:0] _1101;
    wire [3:0] _1104;
    wire [3:0] _1107;
    wire [3:0] _1110;
    wire _1112;
    wire _1113;
    wire _3284;
    wire _3285;
    wire _3286;
    wire _3287;
    wire _129;
    reg _776;
    wire [3:0] _1067;
    wire [3:0] _1064;
    wire [3:0] _1061;
    wire [3:0] _1059;
    wire [3:0] _1062;
    wire [3:0] _1065;
    wire [3:0] _1068;
    wire [3:0] _1071;
    wire [3:0] _1074;
    wire [3:0] _1077;
    wire [3:0] _1080;
    wire _1082;
    wire _1083;
    wire _3288;
    wire _3289;
    wire _3290;
    wire _3291;
    wire _130;
    reg _753;
    wire [3:0] _1328;
    wire [3:0] _1325;
    wire [3:0] _1322;
    wire [3:0] _1318;
    wire [3:0] _1323;
    wire [3:0] _1326;
    wire [3:0] _1329;
    wire [3:0] _1332;
    wire _1334;
    wire _1335;
    wire _3292;
    wire _3293;
    wire _3294;
    wire _3295;
    wire _131;
    reg _1039;
    wire [3:0] _1613;
    wire [3:0] _1610;
    wire [3:0] _1607;
    wire [3:0] _1604;
    wire [3:0] _1600;
    wire [3:0] _1605;
    wire [3:0] _1608;
    wire [3:0] _1611;
    wire [3:0] _1614;
    wire _1616;
    wire _1617;
    wire _3296;
    wire _3297;
    wire _3298;
    wire _3299;
    wire _132;
    reg _1321;
    wire [3:0] _1346;
    wire [3:0] _1343;
    wire [3:0] _1341;
    wire [3:0] _1344;
    wire [3:0] _1347;
    wire [3:0] _1350;
    wire [3:0] _1353;
    wire [3:0] _1356;
    wire [3:0] _1359;
    wire [3:0] _1362;
    wire _1364;
    wire _1365;
    wire _3300;
    wire _3301;
    wire _3302;
    wire _3303;
    wire _133;
    reg _1035;
    wire [3:0] _1382;
    wire [3:0] _1379;
    wire [3:0] _1376;
    wire [3:0] _1373;
    wire [3:0] _1371;
    wire [3:0] _1374;
    wire [3:0] _1377;
    wire [3:0] _1380;
    wire [3:0] _1383;
    wire [3:0] _1386;
    wire [3:0] _1389;
    wire [3:0] _1392;
    wire _1394;
    wire _1395;
    wire _3304;
    wire _3305;
    wire _3306;
    wire _3307;
    wire _134;
    reg _1058;
    wire [3:0] _1412;
    wire [3:0] _1409;
    wire [3:0] _1406;
    wire [3:0] _1403;
    wire [3:0] _1401;
    wire [3:0] _1404;
    wire [3:0] _1407;
    wire [3:0] _1410;
    wire [3:0] _1413;
    wire [3:0] _1416;
    wire [3:0] _1419;
    wire [3:0] _1422;
    wire _1424;
    wire _1425;
    wire _3308;
    wire _3309;
    wire _3310;
    wire _3311;
    wire _135;
    reg _1088;
    wire [3:0] _1442;
    wire [3:0] _1439;
    wire [3:0] _1436;
    wire [3:0] _1433;
    wire [3:0] _1431;
    wire [3:0] _1434;
    wire [3:0] _1437;
    wire [3:0] _1440;
    wire [3:0] _1443;
    wire [3:0] _1446;
    wire [3:0] _1449;
    wire [3:0] _1452;
    wire _1454;
    wire _1455;
    wire _3312;
    wire _3313;
    wire _3314;
    wire _3315;
    wire _136;
    reg _1118;
    wire [3:0] _1472;
    wire [3:0] _1469;
    wire [3:0] _1466;
    wire [3:0] _1463;
    wire [3:0] _1461;
    wire [3:0] _1464;
    wire [3:0] _1467;
    wire [3:0] _1470;
    wire [3:0] _1473;
    wire [3:0] _1476;
    wire [3:0] _1479;
    wire [3:0] _1482;
    wire _1484;
    wire _1485;
    wire _3316;
    wire _3317;
    wire _3318;
    wire _3319;
    wire _137;
    reg _1148;
    wire [3:0] _1502;
    wire [3:0] _1499;
    wire [3:0] _1496;
    wire [3:0] _1493;
    wire [3:0] _1491;
    wire [3:0] _1494;
    wire [3:0] _1497;
    wire [3:0] _1500;
    wire [3:0] _1503;
    wire [3:0] _1506;
    wire [3:0] _1509;
    wire [3:0] _1512;
    wire _1514;
    wire _1515;
    wire _3320;
    wire _3321;
    wire _3322;
    wire _3323;
    wire _138;
    reg _1178;
    wire [3:0] _1532;
    wire [3:0] _1529;
    wire [3:0] _1526;
    wire [3:0] _1523;
    wire [3:0] _1521;
    wire [3:0] _1524;
    wire [3:0] _1527;
    wire [3:0] _1530;
    wire [3:0] _1533;
    wire [3:0] _1536;
    wire [3:0] _1539;
    wire [3:0] _1542;
    wire _1544;
    wire _1545;
    wire _3324;
    wire _3325;
    wire _3326;
    wire _3327;
    wire _139;
    reg _1208;
    wire [3:0] _1562;
    wire [3:0] _1559;
    wire [3:0] _1556;
    wire [3:0] _1553;
    wire [3:0] _1551;
    wire [3:0] _1554;
    wire [3:0] _1557;
    wire [3:0] _1560;
    wire [3:0] _1563;
    wire [3:0] _1566;
    wire [3:0] _1569;
    wire [3:0] _1572;
    wire _1574;
    wire _1575;
    wire _3328;
    wire _3329;
    wire _3330;
    wire _3331;
    wire _140;
    reg _1238;
    wire [3:0] _1584;
    wire [3:0] _1581;
    wire [3:0] _1579;
    wire [3:0] _1582;
    wire [3:0] _1585;
    wire [3:0] _1588;
    wire [3:0] _1591;
    wire _1593;
    wire _1594;
    wire _3332;
    wire _3333;
    wire _3334;
    wire _3335;
    wire _141;
    reg _1268;
    wire [3:0] _1869;
    wire [3:0] _1866;
    wire [3:0] _1863;
    wire [3:0] _1861;
    wire [3:0] _1864;
    wire [3:0] _1867;
    wire [3:0] _1870;
    wire [3:0] _1873;
    wire _1875;
    wire _1876;
    wire _3336;
    wire _3337;
    wire _3338;
    wire _3339;
    wire _142;
    reg _1550;
    wire [3:0] _1841;
    wire [3:0] _1838;
    wire [3:0] _1835;
    wire [3:0] _1833;
    wire [3:0] _1836;
    wire [3:0] _1839;
    wire [3:0] _1842;
    wire [3:0] _1845;
    wire [3:0] _1848;
    wire [3:0] _1851;
    wire [3:0] _1854;
    wire _1856;
    wire _1857;
    wire _3340;
    wire _3341;
    wire _3342;
    wire _3343;
    wire _143;
    reg _1520;
    wire [3:0] _1811;
    wire [3:0] _1808;
    wire [3:0] _1805;
    wire [3:0] _1803;
    wire [3:0] _1806;
    wire [3:0] _1809;
    wire [3:0] _1812;
    wire [3:0] _1815;
    wire [3:0] _1818;
    wire [3:0] _1821;
    wire [3:0] _1824;
    wire _1826;
    wire _1827;
    wire _3344;
    wire _3345;
    wire _3346;
    wire _3347;
    wire _144;
    reg _1490;
    wire [3:0] _1781;
    wire [3:0] _1778;
    wire [3:0] _1775;
    wire [3:0] _1773;
    wire [3:0] _1776;
    wire [3:0] _1779;
    wire [3:0] _1782;
    wire [3:0] _1785;
    wire [3:0] _1788;
    wire [3:0] _1791;
    wire [3:0] _1794;
    wire _1796;
    wire _1797;
    wire _3348;
    wire _3349;
    wire _3350;
    wire _3351;
    wire _145;
    reg _1460;
    wire [3:0] _1751;
    wire [3:0] _1748;
    wire [3:0] _1745;
    wire [3:0] _1743;
    wire [3:0] _1746;
    wire [3:0] _1749;
    wire [3:0] _1752;
    wire [3:0] _1755;
    wire [3:0] _1758;
    wire [3:0] _1761;
    wire [3:0] _1764;
    wire _1766;
    wire _1767;
    wire _3352;
    wire _3353;
    wire _3354;
    wire _3355;
    wire _146;
    reg _1430;
    wire [3:0] _1721;
    wire [3:0] _1718;
    wire [3:0] _1715;
    wire [3:0] _1713;
    wire [3:0] _1716;
    wire [3:0] _1719;
    wire [3:0] _1722;
    wire [3:0] _1725;
    wire [3:0] _1728;
    wire [3:0] _1731;
    wire [3:0] _1734;
    wire _1736;
    wire _1737;
    wire _3356;
    wire _3357;
    wire _3358;
    wire _3359;
    wire _147;
    reg _1400;
    wire [3:0] _1691;
    wire [3:0] _1688;
    wire [3:0] _1685;
    wire [3:0] _1683;
    wire [3:0] _1686;
    wire [3:0] _1689;
    wire [3:0] _1692;
    wire [3:0] _1695;
    wire [3:0] _1698;
    wire [3:0] _1701;
    wire [3:0] _1704;
    wire _1706;
    wire _1707;
    wire _3360;
    wire _3361;
    wire _3362;
    wire _3363;
    wire _148;
    reg _1370;
    wire [3:0] _1661;
    wire [3:0] _1658;
    wire [3:0] _1655;
    wire [3:0] _1653;
    wire [3:0] _1656;
    wire [3:0] _1659;
    wire [3:0] _1662;
    wire [3:0] _1665;
    wire [3:0] _1668;
    wire [3:0] _1671;
    wire [3:0] _1674;
    wire _1676;
    wire _1677;
    wire _3364;
    wire _3365;
    wire _3366;
    wire _3367;
    wire _149;
    reg _1340;
    wire [3:0] _1631;
    wire [3:0] _1628;
    wire [3:0] _1625;
    wire [3:0] _1623;
    wire [3:0] _1626;
    wire [3:0] _1629;
    wire [3:0] _1632;
    wire [3:0] _1635;
    wire [3:0] _1638;
    wire [3:0] _1641;
    wire [3:0] _1644;
    wire _1646;
    wire _1647;
    wire _3368;
    wire _3369;
    wire _3370;
    wire _3371;
    wire _150;
    reg _1317;
    wire [3:0] _1892;
    wire [3:0] _1889;
    wire [3:0] _1886;
    wire [3:0] _1882;
    wire [3:0] _1887;
    wire [3:0] _1890;
    wire [3:0] _1893;
    wire [3:0] _1896;
    wire _1898;
    wire _1899;
    wire _3372;
    wire _3373;
    wire _3374;
    wire _3375;
    wire _151;
    reg _1603;
    wire [3:0] _2177;
    wire [3:0] _2174;
    wire [3:0] _2171;
    wire [3:0] _2168;
    wire [3:0] _2164;
    wire [3:0] _2169;
    wire [3:0] _2172;
    wire [3:0] _2175;
    wire [3:0] _2178;
    wire _2180;
    wire _2181;
    wire _3376;
    wire _3377;
    wire _3378;
    wire _3379;
    wire _152;
    reg _1885;
    wire [3:0] _1910;
    wire [3:0] _1907;
    wire [3:0] _1905;
    wire [3:0] _1908;
    wire [3:0] _1911;
    wire [3:0] _1914;
    wire [3:0] _1917;
    wire [3:0] _1920;
    wire [3:0] _1923;
    wire [3:0] _1926;
    wire _1928;
    wire _1929;
    wire _3380;
    wire _3381;
    wire _3382;
    wire _3383;
    wire _153;
    reg _1599;
    wire [3:0] _1946;
    wire [3:0] _1943;
    wire [3:0] _1940;
    wire [3:0] _1937;
    wire [3:0] _1935;
    wire [3:0] _1938;
    wire [3:0] _1941;
    wire [3:0] _1944;
    wire [3:0] _1947;
    wire [3:0] _1950;
    wire [3:0] _1953;
    wire [3:0] _1956;
    wire _1958;
    wire _1959;
    wire _3384;
    wire _3385;
    wire _3386;
    wire _3387;
    wire _154;
    reg _1622;
    wire [3:0] _1976;
    wire [3:0] _1973;
    wire [3:0] _1970;
    wire [3:0] _1967;
    wire [3:0] _1965;
    wire [3:0] _1968;
    wire [3:0] _1971;
    wire [3:0] _1974;
    wire [3:0] _1977;
    wire [3:0] _1980;
    wire [3:0] _1983;
    wire [3:0] _1986;
    wire _1988;
    wire _1989;
    wire _3388;
    wire _3389;
    wire _3390;
    wire _3391;
    wire _155;
    reg _1652;
    wire [3:0] _2006;
    wire [3:0] _2003;
    wire [3:0] _2000;
    wire [3:0] _1997;
    wire [3:0] _1995;
    wire [3:0] _1998;
    wire [3:0] _2001;
    wire [3:0] _2004;
    wire [3:0] _2007;
    wire [3:0] _2010;
    wire [3:0] _2013;
    wire [3:0] _2016;
    wire _2018;
    wire _2019;
    wire _3392;
    wire _3393;
    wire _3394;
    wire _3395;
    wire _156;
    reg _1682;
    wire [3:0] _2036;
    wire [3:0] _2033;
    wire [3:0] _2030;
    wire [3:0] _2027;
    wire [3:0] _2025;
    wire [3:0] _2028;
    wire [3:0] _2031;
    wire [3:0] _2034;
    wire [3:0] _2037;
    wire [3:0] _2040;
    wire [3:0] _2043;
    wire [3:0] _2046;
    wire _2048;
    wire _2049;
    wire _3396;
    wire _3397;
    wire _3398;
    wire _3399;
    wire _157;
    reg _1712;
    wire [3:0] _2066;
    wire [3:0] _2063;
    wire [3:0] _2060;
    wire [3:0] _2057;
    wire [3:0] _2055;
    wire [3:0] _2058;
    wire [3:0] _2061;
    wire [3:0] _2064;
    wire [3:0] _2067;
    wire [3:0] _2070;
    wire [3:0] _2073;
    wire [3:0] _2076;
    wire _2078;
    wire _2079;
    wire _3400;
    wire _3401;
    wire _3402;
    wire _3403;
    wire _158;
    reg _1742;
    wire [3:0] _2096;
    wire [3:0] _2093;
    wire [3:0] _2090;
    wire [3:0] _2087;
    wire [3:0] _2085;
    wire [3:0] _2088;
    wire [3:0] _2091;
    wire [3:0] _2094;
    wire [3:0] _2097;
    wire [3:0] _2100;
    wire [3:0] _2103;
    wire [3:0] _2106;
    wire _2108;
    wire _2109;
    wire _3404;
    wire _3405;
    wire _3406;
    wire _3407;
    wire _159;
    reg _1772;
    wire [3:0] _2126;
    wire [3:0] _2123;
    wire [3:0] _2120;
    wire [3:0] _2117;
    wire [3:0] _2115;
    wire [3:0] _2118;
    wire [3:0] _2121;
    wire [3:0] _2124;
    wire [3:0] _2127;
    wire [3:0] _2130;
    wire [3:0] _2133;
    wire [3:0] _2136;
    wire _2138;
    wire _2139;
    wire _3408;
    wire _3409;
    wire _3410;
    wire _3411;
    wire _160;
    reg _1802;
    wire [3:0] _2148;
    wire [3:0] _2145;
    wire [3:0] _2143;
    wire [3:0] _2146;
    wire [3:0] _2149;
    wire [3:0] _2152;
    wire [3:0] _2155;
    wire _2157;
    wire _2158;
    wire _3412;
    wire _3413;
    wire _3414;
    wire _3415;
    wire _161;
    reg _1832;
    wire [3:0] _2433;
    wire [3:0] _2430;
    wire [3:0] _2427;
    wire [3:0] _2425;
    wire [3:0] _2428;
    wire [3:0] _2431;
    wire [3:0] _2434;
    wire [3:0] _2437;
    wire _2439;
    wire _2440;
    wire _3416;
    wire _3417;
    wire _3418;
    wire _3419;
    wire _162;
    reg _2114;
    wire [3:0] _2405;
    wire [3:0] _2402;
    wire [3:0] _2399;
    wire [3:0] _2397;
    wire [3:0] _2400;
    wire [3:0] _2403;
    wire [3:0] _2406;
    wire [3:0] _2409;
    wire [3:0] _2412;
    wire [3:0] _2415;
    wire [3:0] _2418;
    wire _2420;
    wire _2421;
    wire _3420;
    wire _3421;
    wire _3422;
    wire _3423;
    wire _163;
    reg _2084;
    wire [3:0] _2375;
    wire [3:0] _2372;
    wire [3:0] _2369;
    wire [3:0] _2367;
    wire [3:0] _2370;
    wire [3:0] _2373;
    wire [3:0] _2376;
    wire [3:0] _2379;
    wire [3:0] _2382;
    wire [3:0] _2385;
    wire [3:0] _2388;
    wire _2390;
    wire _2391;
    wire _3424;
    wire _3425;
    wire _3426;
    wire _3427;
    wire _164;
    reg _2054;
    wire [3:0] _2345;
    wire [3:0] _2342;
    wire [3:0] _2339;
    wire [3:0] _2337;
    wire [3:0] _2340;
    wire [3:0] _2343;
    wire [3:0] _2346;
    wire [3:0] _2349;
    wire [3:0] _2352;
    wire [3:0] _2355;
    wire [3:0] _2358;
    wire _2360;
    wire _2361;
    wire _3428;
    wire _3429;
    wire _3430;
    wire _3431;
    wire _165;
    reg _2024;
    wire [3:0] _2315;
    wire [3:0] _2312;
    wire [3:0] _2309;
    wire [3:0] _2307;
    wire [3:0] _2310;
    wire [3:0] _2313;
    wire [3:0] _2316;
    wire [3:0] _2319;
    wire [3:0] _2322;
    wire [3:0] _2325;
    wire [3:0] _2328;
    wire _2330;
    wire _2331;
    wire _3432;
    wire _3433;
    wire _3434;
    wire _3435;
    wire _166;
    reg _1994;
    wire [3:0] _2285;
    wire [3:0] _2282;
    wire [3:0] _2279;
    wire [3:0] _2277;
    wire [3:0] _2280;
    wire [3:0] _2283;
    wire [3:0] _2286;
    wire [3:0] _2289;
    wire [3:0] _2292;
    wire [3:0] _2295;
    wire [3:0] _2298;
    wire _2300;
    wire _2301;
    wire _3436;
    wire _3437;
    wire _3438;
    wire _3439;
    wire _167;
    reg _1964;
    wire [3:0] _2255;
    wire [3:0] _2252;
    wire [3:0] _2249;
    wire [3:0] _2247;
    wire [3:0] _2250;
    wire [3:0] _2253;
    wire [3:0] _2256;
    wire [3:0] _2259;
    wire [3:0] _2262;
    wire [3:0] _2265;
    wire [3:0] _2268;
    wire _2270;
    wire _2271;
    wire _3440;
    wire _3441;
    wire _3442;
    wire _3443;
    wire _168;
    reg _1934;
    wire [3:0] _2225;
    wire [3:0] _2222;
    wire [3:0] _2219;
    wire [3:0] _2217;
    wire [3:0] _2220;
    wire [3:0] _2223;
    wire [3:0] _2226;
    wire [3:0] _2229;
    wire [3:0] _2232;
    wire [3:0] _2235;
    wire [3:0] _2238;
    wire _2240;
    wire _2241;
    wire _3444;
    wire _3445;
    wire _3446;
    wire _3447;
    wire _169;
    reg _1904;
    wire [3:0] _2195;
    wire [3:0] _2192;
    wire [3:0] _2189;
    wire [3:0] _2187;
    wire [3:0] _2190;
    wire [3:0] _2193;
    wire [3:0] _2196;
    wire [3:0] _2199;
    wire [3:0] _2202;
    wire [3:0] _2205;
    wire [3:0] _2208;
    wire _2210;
    wire _2211;
    wire _3448;
    wire _3449;
    wire _3450;
    wire _3451;
    wire _170;
    reg _1881;
    wire [3:0] _2456;
    wire [3:0] _2453;
    wire [3:0] _2450;
    wire [3:0] _2446;
    wire [3:0] _2451;
    wire [3:0] _2454;
    wire [3:0] _2457;
    wire [3:0] _2460;
    wire _2462;
    wire _2463;
    wire _3452;
    wire _3453;
    wire _3454;
    wire _3455;
    wire _171;
    reg _2167;
    wire [3:0] _2741;
    wire [3:0] _2738;
    wire [3:0] _2735;
    wire [3:0] _2732;
    wire [3:0] _2728;
    wire [3:0] _2733;
    wire [3:0] _2736;
    wire [3:0] _2739;
    wire [3:0] _2742;
    wire _2744;
    wire _2745;
    wire _3456;
    wire _3457;
    wire _3458;
    wire _3459;
    wire _172;
    reg _2449;
    wire [3:0] _2474;
    wire [3:0] _2471;
    wire [3:0] _2469;
    wire [3:0] _2472;
    wire [3:0] _2475;
    wire [3:0] _2478;
    wire [3:0] _2481;
    wire [3:0] _2484;
    wire [3:0] _2487;
    wire [3:0] _2490;
    wire _2492;
    wire _2493;
    wire _3460;
    wire _3461;
    wire _3462;
    wire _3463;
    wire _173;
    reg _2163;
    wire [3:0] _2510;
    wire [3:0] _2507;
    wire [3:0] _2504;
    wire [3:0] _2501;
    wire [3:0] _2499;
    wire [3:0] _2502;
    wire [3:0] _2505;
    wire [3:0] _2508;
    wire [3:0] _2511;
    wire [3:0] _2514;
    wire [3:0] _2517;
    wire [3:0] _2520;
    wire _2522;
    wire _2523;
    wire _3464;
    wire _3465;
    wire _3466;
    wire _3467;
    wire _174;
    reg _2186;
    wire [3:0] _2540;
    wire [3:0] _2537;
    wire [3:0] _2534;
    wire [3:0] _2531;
    wire [3:0] _2529;
    wire [3:0] _2532;
    wire [3:0] _2535;
    wire [3:0] _2538;
    wire [3:0] _2541;
    wire [3:0] _2544;
    wire [3:0] _2547;
    wire [3:0] _2550;
    wire _2552;
    wire _2553;
    wire _3468;
    wire _3469;
    wire _3470;
    wire _3471;
    wire _175;
    reg _2216;
    wire [3:0] _2570;
    wire [3:0] _2567;
    wire [3:0] _2564;
    wire [3:0] _2561;
    wire [3:0] _2559;
    wire [3:0] _2562;
    wire [3:0] _2565;
    wire [3:0] _2568;
    wire [3:0] _2571;
    wire [3:0] _2574;
    wire [3:0] _2577;
    wire [3:0] _2580;
    wire _2582;
    wire _2583;
    wire _3472;
    wire _3473;
    wire _3474;
    wire _3475;
    wire _176;
    reg _2246;
    wire [3:0] _2600;
    wire [3:0] _2597;
    wire [3:0] _2594;
    wire [3:0] _2591;
    wire [3:0] _2589;
    wire [3:0] _2592;
    wire [3:0] _2595;
    wire [3:0] _2598;
    wire [3:0] _2601;
    wire [3:0] _2604;
    wire [3:0] _2607;
    wire [3:0] _2610;
    wire _2612;
    wire _2613;
    wire _3476;
    wire _3477;
    wire _3478;
    wire _3479;
    wire _177;
    reg _2276;
    wire [3:0] _2630;
    wire [3:0] _2627;
    wire [3:0] _2624;
    wire [3:0] _2621;
    wire [3:0] _2619;
    wire [3:0] _2622;
    wire [3:0] _2625;
    wire [3:0] _2628;
    wire [3:0] _2631;
    wire [3:0] _2634;
    wire [3:0] _2637;
    wire [3:0] _2640;
    wire _2642;
    wire _2643;
    wire _3480;
    wire _3481;
    wire _3482;
    wire _3483;
    wire _178;
    reg _2306;
    wire [3:0] _2660;
    wire [3:0] _2657;
    wire [3:0] _2654;
    wire [3:0] _2651;
    wire [3:0] _2649;
    wire [3:0] _2652;
    wire [3:0] _2655;
    wire [3:0] _2658;
    wire [3:0] _2661;
    wire [3:0] _2664;
    wire [3:0] _2667;
    wire [3:0] _2670;
    wire _2672;
    wire _2673;
    wire _3484;
    wire _3485;
    wire _3486;
    wire _3487;
    wire _179;
    reg _2336;
    wire [3:0] _2690;
    wire [3:0] _2687;
    wire [3:0] _2684;
    wire [3:0] _2681;
    wire [3:0] _2679;
    wire [3:0] _2682;
    wire [3:0] _2685;
    wire [3:0] _2688;
    wire [3:0] _2691;
    wire [3:0] _2694;
    wire [3:0] _2697;
    wire [3:0] _2700;
    wire _2702;
    wire _2703;
    wire _3488;
    wire _3489;
    wire _3490;
    wire _3491;
    wire _180;
    reg _2366;
    wire [3:0] _2712;
    wire [3:0] _2709;
    wire [3:0] _2707;
    wire [3:0] _2710;
    wire [3:0] _2713;
    wire [3:0] _2716;
    wire [3:0] _2719;
    wire _2721;
    wire _2722;
    wire _3492;
    wire _3493;
    wire _3494;
    wire _3495;
    wire _181;
    reg _2396;
    wire [3:0] _2997;
    wire [3:0] _2994;
    wire [3:0] _2991;
    wire [3:0] _2989;
    wire [3:0] _2992;
    wire [3:0] _2995;
    wire [3:0] _2998;
    wire [3:0] _3001;
    wire _3003;
    wire _3004;
    wire _3496;
    wire _3497;
    wire _3498;
    wire _3499;
    wire _182;
    reg _2678;
    wire [3:0] _2969;
    wire [3:0] _2966;
    wire [3:0] _2963;
    wire [3:0] _2961;
    wire [3:0] _2964;
    wire [3:0] _2967;
    wire [3:0] _2970;
    wire [3:0] _2973;
    wire [3:0] _2976;
    wire [3:0] _2979;
    wire [3:0] _2982;
    wire _2984;
    wire _2985;
    wire _3500;
    wire _3501;
    wire _3502;
    wire _3503;
    wire _183;
    reg _2648;
    wire [3:0] _2939;
    wire [3:0] _2936;
    wire [3:0] _2933;
    wire [3:0] _2931;
    wire [3:0] _2934;
    wire [3:0] _2937;
    wire [3:0] _2940;
    wire [3:0] _2943;
    wire [3:0] _2946;
    wire [3:0] _2949;
    wire [3:0] _2952;
    wire _2954;
    wire _2955;
    wire _3504;
    wire _3505;
    wire _3506;
    wire _3507;
    wire _184;
    reg _2618;
    wire [3:0] _2909;
    wire [3:0] _2906;
    wire [3:0] _2903;
    wire [3:0] _2901;
    wire [3:0] _2904;
    wire [3:0] _2907;
    wire [3:0] _2910;
    wire [3:0] _2913;
    wire [3:0] _2916;
    wire [3:0] _2919;
    wire [3:0] _2922;
    wire _2924;
    wire _2925;
    wire _3508;
    wire _3509;
    wire _3510;
    wire _3511;
    wire _185;
    reg _2588;
    wire [3:0] _2879;
    wire [3:0] _2876;
    wire [3:0] _2873;
    wire [3:0] _2871;
    wire [3:0] _2874;
    wire [3:0] _2877;
    wire [3:0] _2880;
    wire [3:0] _2883;
    wire [3:0] _2886;
    wire [3:0] _2889;
    wire [3:0] _2892;
    wire _2894;
    wire _2895;
    wire _3512;
    wire _3513;
    wire _3514;
    wire _3515;
    wire _186;
    reg _2558;
    wire [3:0] _2849;
    wire [3:0] _2846;
    wire [3:0] _2843;
    wire [3:0] _2841;
    wire [3:0] _2844;
    wire [3:0] _2847;
    wire [3:0] _2850;
    wire [3:0] _2853;
    wire [3:0] _2856;
    wire [3:0] _2859;
    wire [3:0] _2862;
    wire _2864;
    wire _2865;
    wire _3516;
    wire _3517;
    wire _3518;
    wire _3519;
    wire _187;
    reg _2528;
    wire [3:0] _2819;
    wire [3:0] _2816;
    wire [3:0] _2813;
    wire [3:0] _2811;
    wire [3:0] _2814;
    wire [3:0] _2817;
    wire [3:0] _2820;
    wire [3:0] _2823;
    wire [3:0] _2826;
    wire [3:0] _2829;
    wire [3:0] _2832;
    wire _2834;
    wire _2835;
    wire _3520;
    wire _3521;
    wire _3522;
    wire _3523;
    wire _188;
    reg _2498;
    wire [3:0] _2789;
    wire [3:0] _2786;
    wire [3:0] _2783;
    wire [3:0] _2781;
    wire [3:0] _2784;
    wire [3:0] _2787;
    wire [3:0] _2790;
    wire [3:0] _2793;
    wire [3:0] _2796;
    wire [3:0] _2799;
    wire [3:0] _2802;
    wire _2804;
    wire _2805;
    wire _3524;
    wire _3525;
    wire _3526;
    wire _3527;
    wire _189;
    reg _2468;
    wire [3:0] _2759;
    wire [3:0] _2756;
    wire [3:0] _2753;
    wire [3:0] _2751;
    wire [3:0] _2754;
    wire [3:0] _2757;
    wire [3:0] _2760;
    wire [3:0] _2763;
    wire [3:0] _2766;
    wire [3:0] _2769;
    wire [3:0] _2772;
    wire _2774;
    wire _2775;
    wire _3528;
    wire _3529;
    wire _3530;
    wire _3531;
    wire _190;
    reg _2445;
    wire [3:0] _3010;
    wire [3:0] _3008;
    wire [3:0] _3011;
    wire [3:0] _3014;
    wire _3016;
    wire _3017;
    wire _3532;
    wire _3533;
    wire _3534;
    wire _3535;
    wire _191;
    reg _2731;
    wire [3:0] _3023;
    wire [3:0] _3021;
    wire [3:0] _3024;
    wire [3:0] _3027;
    wire [3:0] _3030;
    wire [3:0] _3033;
    wire _3035;
    wire _3036;
    wire _3536;
    wire _3537;
    wire _3538;
    wire _3539;
    wire _192;
    reg _2727;
    wire [3:0] _3042;
    wire [3:0] _3040;
    wire [3:0] _3043;
    wire [3:0] _3046;
    wire [3:0] _3049;
    wire [3:0] _3052;
    wire _3054;
    wire _3055;
    wire _3540;
    wire _3541;
    wire _3542;
    wire _3543;
    wire _193;
    reg _2750;
    wire [3:0] _3061;
    wire [3:0] _3059;
    wire [3:0] _3062;
    wire [3:0] _3065;
    wire [3:0] _3068;
    wire [3:0] _3071;
    wire _3073;
    wire _3074;
    wire _3544;
    wire _3545;
    wire _3546;
    wire _3547;
    wire _194;
    reg _2780;
    wire [3:0] _3080;
    wire [3:0] _3078;
    wire [3:0] _3081;
    wire [3:0] _3084;
    wire [3:0] _3087;
    wire [3:0] _3090;
    wire _3092;
    wire _3093;
    wire _3548;
    wire _3549;
    wire _3550;
    wire _3551;
    wire _195;
    reg _2810;
    wire [3:0] _3099;
    wire [3:0] _3097;
    wire [3:0] _3100;
    wire [3:0] _3103;
    wire [3:0] _3106;
    wire [3:0] _3109;
    wire _3111;
    wire _3112;
    wire _3552;
    wire _3553;
    wire _3554;
    wire _3555;
    wire _196;
    reg _2840;
    wire [3:0] _3118;
    wire [3:0] _3116;
    wire [3:0] _3119;
    wire [3:0] _3122;
    wire [3:0] _3125;
    wire [3:0] _3128;
    wire _3130;
    wire _3131;
    wire _3556;
    wire _3557;
    wire _3558;
    wire _3559;
    wire _197;
    reg _2870;
    wire [3:0] _3137;
    wire [3:0] _3135;
    wire [3:0] _3138;
    wire [3:0] _3141;
    wire [3:0] _3144;
    wire [3:0] _3147;
    wire _3149;
    wire _3150;
    wire _3560;
    wire _3561;
    wire _3562;
    wire _3563;
    wire _198;
    reg _2900;
    wire [3:0] _3156;
    wire [3:0] _3154;
    wire [3:0] _3157;
    wire [3:0] _3160;
    wire [3:0] _3163;
    wire [3:0] _3166;
    wire _3168;
    wire _3169;
    wire _3564;
    wire _3565;
    wire _3566;
    wire _3567;
    wire _199;
    reg _2930;
    wire [3:0] _3569;
    wire [3:0] _3572;
    wire [3:0] _3575;
    wire _3577;
    wire _222;
    wire _223;
    wire _3582;
    wire _3579;
    wire _3580;
    wire _3581;
    wire _3583;
    wire _200;
    reg _2960;
    wire _3578;
    wire gnd;
    wire _3584;
    wire [3:0] _529;
    wire _530;
    wire _531;
    wire _3585;
    wire _201;
    wire [15:0] _229;
    wire [15:0] _232;
    wire [15:0] _235;
    wire [15:0] _238;
    wire [15:0] _241;
    wire [15:0] _244;
    wire [15:0] _247;
    wire [15:0] _250;
    wire [15:0] _253;
    wire [15:0] _256;
    wire [15:0] _259;
    wire [15:0] _262;
    wire [15:0] _265;
    wire [15:0] _268;
    wire [15:0] _271;
    wire [15:0] _274;
    wire [15:0] _277;
    wire [15:0] _280;
    wire [15:0] _283;
    wire [15:0] _286;
    wire [15:0] _289;
    wire [15:0] _292;
    wire [15:0] _295;
    wire [15:0] _298;
    wire [15:0] _301;
    wire [15:0] _304;
    wire [15:0] _307;
    wire [15:0] _310;
    wire [15:0] _313;
    wire [15:0] _316;
    wire [15:0] _319;
    wire [15:0] _322;
    wire [15:0] _325;
    wire [15:0] _328;
    wire [15:0] _331;
    wire [15:0] _334;
    wire [15:0] _337;
    wire [15:0] _340;
    wire [15:0] _343;
    wire [15:0] _346;
    wire [15:0] _349;
    wire [15:0] _352;
    wire [15:0] _355;
    wire [15:0] _358;
    wire [15:0] _361;
    wire [15:0] _364;
    wire [15:0] _367;
    wire [15:0] _370;
    wire [15:0] _373;
    wire [15:0] _376;
    wire [15:0] _379;
    wire [15:0] _382;
    wire [15:0] _385;
    wire [15:0] _388;
    wire [15:0] _391;
    wire [15:0] _394;
    wire [15:0] _397;
    wire [15:0] _400;
    wire [15:0] _403;
    wire [15:0] _406;
    wire [15:0] _409;
    wire [15:0] _412;
    wire [15:0] _415;
    wire [15:0] _418;
    wire [15:0] _421;
    wire [15:0] _424;
    wire [15:0] _427;
    wire [15:0] _430;
    wire [15:0] _433;
    wire [15:0] _436;
    wire [15:0] _439;
    wire [15:0] _442;
    wire [15:0] _445;
    wire [15:0] _448;
    wire [15:0] _451;
    wire [15:0] _454;
    wire [15:0] _457;
    wire [15:0] _460;
    wire [15:0] _463;
    wire [15:0] _466;
    wire [15:0] _469;
    wire [15:0] _472;
    wire [15:0] _475;
    wire [15:0] _478;
    wire [15:0] _481;
    wire [15:0] _484;
    wire [15:0] _487;
    wire [15:0] _490;
    wire [15:0] _493;
    wire [15:0] _496;
    wire [15:0] _499;
    wire [15:0] _502;
    wire [15:0] _505;
    wire [15:0] _508;
    wire [15:0] _511;
    wire [15:0] _514;
    wire [15:0] _517;
    wire [15:0] _520;
    wire [15:0] _523;
    wire [15:0] _526;
    wire _3589;
    wire _221;
    wire _3590;
    wire [30:0] _3587;
    wire [31:0] _3591;
    wire [31:0] _3586;
    wire [3:0] _217;
    wire [3:0] _203;
    wire _218;
    wire _205;
    wire _219;
    wire _207;
    wire _209;
    wire [31:0] _211;
    wire [31:0] _212;
    reg [31:0] _220;
    wire [3:0] _214;
    reg [31:0] _3895;
    assign _3891 = 15'b000000000000000;
    assign _3892 = { _3891,
                     _534 };
    assign _3889 = { _3891,
                     _546 };
    assign _3886 = { _3891,
                     _566 };
    assign _3883 = { _3891,
                     _589 };
    assign _3880 = { _3891,
                     _612 };
    assign _3877 = { _3891,
                     _635 };
    assign _3874 = { _3891,
                     _658 };
    assign _3871 = { _3891,
                     _681 };
    assign _3868 = { _3891,
                     _704 };
    assign _3865 = { _3891,
                     _727 };
    assign _3862 = { _3891,
                     _541 };
    assign _3859 = { _3891,
                     _537 };
    assign _3856 = { _3891,
                     _556 };
    assign _3853 = { _3891,
                     _579 };
    assign _3850 = { _3891,
                     _602 };
    assign _3847 = { _3891,
                     _625 };
    assign _3844 = { _3891,
                     _648 };
    assign _3841 = { _3891,
                     _671 };
    assign _3838 = { _3891,
                     _694 };
    assign _3835 = { _3891,
                     _717 };
    assign _3832 = { _3891,
                     _757 };
    assign _3829 = { _3891,
                     _753 };
    assign _3826 = { _3891,
                     _776 };
    assign _3823 = { _3891,
                     _806 };
    assign _3820 = { _3891,
                     _836 };
    assign _3817 = { _3891,
                     _866 };
    assign _3814 = { _3891,
                     _896 };
    assign _3811 = { _3891,
                     _926 };
    assign _3808 = { _3891,
                     _956 };
    assign _3805 = { _3891,
                     _986 };
    assign _3802 = { _3891,
                     _1039 };
    assign _3799 = { _3891,
                     _1035 };
    assign _3796 = { _3891,
                     _1058 };
    assign _3793 = { _3891,
                     _1088 };
    assign _3790 = { _3891,
                     _1118 };
    assign _3787 = { _3891,
                     _1148 };
    assign _3784 = { _3891,
                     _1178 };
    assign _3781 = { _3891,
                     _1208 };
    assign _3778 = { _3891,
                     _1238 };
    assign _3775 = { _3891,
                     _1268 };
    assign _3772 = { _3891,
                     _1321 };
    assign _3769 = { _3891,
                     _1317 };
    assign _3766 = { _3891,
                     _1340 };
    assign _3763 = { _3891,
                     _1370 };
    assign _3760 = { _3891,
                     _1400 };
    assign _3757 = { _3891,
                     _1430 };
    assign _3754 = { _3891,
                     _1460 };
    assign _3751 = { _3891,
                     _1490 };
    assign _3748 = { _3891,
                     _1520 };
    assign _3745 = { _3891,
                     _1550 };
    assign _3742 = { _3891,
                     _1603 };
    assign _3739 = { _3891,
                     _1599 };
    assign _3736 = { _3891,
                     _1622 };
    assign _3733 = { _3891,
                     _1652 };
    assign _3730 = { _3891,
                     _1682 };
    assign _3727 = { _3891,
                     _1712 };
    assign _3724 = { _3891,
                     _1742 };
    assign _3721 = { _3891,
                     _1772 };
    assign _3718 = { _3891,
                     _1802 };
    assign _3715 = { _3891,
                     _1832 };
    assign _3712 = { _3891,
                     _1885 };
    assign _3709 = { _3891,
                     _1881 };
    assign _3706 = { _3891,
                     _1904 };
    assign _3703 = { _3891,
                     _1934 };
    assign _3700 = { _3891,
                     _1964 };
    assign _3697 = { _3891,
                     _1994 };
    assign _3694 = { _3891,
                     _2024 };
    assign _3691 = { _3891,
                     _2054 };
    assign _3688 = { _3891,
                     _2084 };
    assign _3685 = { _3891,
                     _2114 };
    assign _3682 = { _3891,
                     _2167 };
    assign _3679 = { _3891,
                     _2163 };
    assign _3676 = { _3891,
                     _2186 };
    assign _3673 = { _3891,
                     _2216 };
    assign _3670 = { _3891,
                     _2246 };
    assign _3667 = { _3891,
                     _2276 };
    assign _3664 = { _3891,
                     _2306 };
    assign _3661 = { _3891,
                     _2336 };
    assign _3658 = { _3891,
                     _2366 };
    assign _3655 = { _3891,
                     _2396 };
    assign _3652 = { _3891,
                     _2449 };
    assign _3649 = { _3891,
                     _2445 };
    assign _3646 = { _3891,
                     _2468 };
    assign _3643 = { _3891,
                     _2498 };
    assign _3640 = { _3891,
                     _2528 };
    assign _3637 = { _3891,
                     _2558 };
    assign _3634 = { _3891,
                     _2588 };
    assign _3631 = { _3891,
                     _2618 };
    assign _3628 = { _3891,
                     _2648 };
    assign _3625 = { _3891,
                     _2678 };
    assign _3622 = { _3891,
                     _2731 };
    assign _3619 = { _3891,
                     _2727 };
    assign _3616 = { _3891,
                     _2750 };
    assign _3613 = { _3891,
                     _2780 };
    assign _3610 = { _3891,
                     _2810 };
    assign _3607 = { _3891,
                     _2840 };
    assign _3604 = { _3891,
                     _2870 };
    assign _3601 = { _3891,
                     _2900 };
    assign _3598 = { _3891,
                     _2930 };
    assign _3596 = { _3891,
                     _2960 };
    assign _3599 = _3596 + _3598;
    assign _3602 = _3599 + _3601;
    assign _3605 = _3602 + _3604;
    assign _3608 = _3605 + _3607;
    assign _3611 = _3608 + _3610;
    assign _3614 = _3611 + _3613;
    assign _3617 = _3614 + _3616;
    assign _3620 = _3617 + _3619;
    assign _3623 = _3620 + _3622;
    assign _3626 = _3623 + _3625;
    assign _3629 = _3626 + _3628;
    assign _3632 = _3629 + _3631;
    assign _3635 = _3632 + _3634;
    assign _3638 = _3635 + _3637;
    assign _3641 = _3638 + _3640;
    assign _3644 = _3641 + _3643;
    assign _3647 = _3644 + _3646;
    assign _3650 = _3647 + _3649;
    assign _3653 = _3650 + _3652;
    assign _3656 = _3653 + _3655;
    assign _3659 = _3656 + _3658;
    assign _3662 = _3659 + _3661;
    assign _3665 = _3662 + _3664;
    assign _3668 = _3665 + _3667;
    assign _3671 = _3668 + _3670;
    assign _3674 = _3671 + _3673;
    assign _3677 = _3674 + _3676;
    assign _3680 = _3677 + _3679;
    assign _3683 = _3680 + _3682;
    assign _3686 = _3683 + _3685;
    assign _3689 = _3686 + _3688;
    assign _3692 = _3689 + _3691;
    assign _3695 = _3692 + _3694;
    assign _3698 = _3695 + _3697;
    assign _3701 = _3698 + _3700;
    assign _3704 = _3701 + _3703;
    assign _3707 = _3704 + _3706;
    assign _3710 = _3707 + _3709;
    assign _3713 = _3710 + _3712;
    assign _3716 = _3713 + _3715;
    assign _3719 = _3716 + _3718;
    assign _3722 = _3719 + _3721;
    assign _3725 = _3722 + _3724;
    assign _3728 = _3725 + _3727;
    assign _3731 = _3728 + _3730;
    assign _3734 = _3731 + _3733;
    assign _3737 = _3734 + _3736;
    assign _3740 = _3737 + _3739;
    assign _3743 = _3740 + _3742;
    assign _3746 = _3743 + _3745;
    assign _3749 = _3746 + _3748;
    assign _3752 = _3749 + _3751;
    assign _3755 = _3752 + _3754;
    assign _3758 = _3755 + _3757;
    assign _3761 = _3758 + _3760;
    assign _3764 = _3761 + _3763;
    assign _3767 = _3764 + _3766;
    assign _3770 = _3767 + _3769;
    assign _3773 = _3770 + _3772;
    assign _3776 = _3773 + _3775;
    assign _3779 = _3776 + _3778;
    assign _3782 = _3779 + _3781;
    assign _3785 = _3782 + _3784;
    assign _3788 = _3785 + _3787;
    assign _3791 = _3788 + _3790;
    assign _3794 = _3791 + _3793;
    assign _3797 = _3794 + _3796;
    assign _3800 = _3797 + _3799;
    assign _3803 = _3800 + _3802;
    assign _3806 = _3803 + _3805;
    assign _3809 = _3806 + _3808;
    assign _3812 = _3809 + _3811;
    assign _3815 = _3812 + _3814;
    assign _3818 = _3815 + _3817;
    assign _3821 = _3818 + _3820;
    assign _3824 = _3821 + _3823;
    assign _3827 = _3824 + _3826;
    assign _3830 = _3827 + _3829;
    assign _3833 = _3830 + _3832;
    assign _3836 = _3833 + _3835;
    assign _3839 = _3836 + _3838;
    assign _3842 = _3839 + _3841;
    assign _3845 = _3842 + _3844;
    assign _3848 = _3845 + _3847;
    assign _3851 = _3848 + _3850;
    assign _3854 = _3851 + _3853;
    assign _3857 = _3854 + _3856;
    assign _3860 = _3857 + _3859;
    assign _3863 = _3860 + _3862;
    assign _3866 = _3863 + _3865;
    assign _3869 = _3866 + _3868;
    assign _3872 = _3869 + _3871;
    assign _3875 = _3872 + _3874;
    assign _3878 = _3875 + _3877;
    assign _3881 = _3878 + _3880;
    assign _3884 = _3881 + _3883;
    assign _3887 = _3884 + _3886;
    assign _3890 = _3887 + _3889;
    assign _3893 = _3890 + _3892;
    assign _3594 = 16'b0000000000000000;
    assign _3894 = { _3594,
                     _3893 };
    assign _527 = _225 + _526;
    assign _227 = _223 ? _3594 : _225;
    assign _528 = _221 ? _527 : _227;
    assign _1 = _528;
    always @(posedge _209) begin
        if (_223)
            _225 <= _3594;
        else
            _225 <= _1;
    end
    assign _3593 = { _3594,
                     _225 };
    assign _552 = _221 ? _551 : gnd;
    assign _553 = _531 ? gnd : _552;
    assign _2 = _553;
    assign _525 = { _3891,
                    _2 };
    assign _575 = _221 ? _574 : gnd;
    assign _576 = _531 ? gnd : _575;
    assign _3 = _576;
    assign _522 = { _3891,
                    _3 };
    assign _598 = _221 ? _597 : gnd;
    assign _599 = _531 ? gnd : _598;
    assign _4 = _599;
    assign _519 = { _3891,
                    _4 };
    assign _621 = _221 ? _620 : gnd;
    assign _622 = _531 ? gnd : _621;
    assign _5 = _622;
    assign _516 = { _3891,
                    _5 };
    assign _644 = _221 ? _643 : gnd;
    assign _645 = _531 ? gnd : _644;
    assign _6 = _645;
    assign _513 = { _3891,
                    _6 };
    assign _667 = _221 ? _666 : gnd;
    assign _668 = _531 ? gnd : _667;
    assign _7 = _668;
    assign _510 = { _3891,
                    _7 };
    assign _690 = _221 ? _689 : gnd;
    assign _691 = _531 ? gnd : _690;
    assign _8 = _691;
    assign _507 = { _3891,
                    _8 };
    assign _713 = _221 ? _712 : gnd;
    assign _714 = _531 ? gnd : _713;
    assign _9 = _714;
    assign _504 = { _3891,
                    _9 };
    assign _736 = _221 ? _735 : gnd;
    assign _737 = _531 ? gnd : _736;
    assign _10 = _737;
    assign _501 = { _3891,
                    _10 };
    assign _749 = _221 ? _748 : gnd;
    assign _750 = _531 ? gnd : _749;
    assign _11 = _750;
    assign _498 = { _3891,
                    _11 };
    assign _772 = _221 ? _771 : gnd;
    assign _773 = _531 ? gnd : _772;
    assign _12 = _773;
    assign _495 = { _3891,
                    _12 };
    assign _802 = _221 ? _801 : gnd;
    assign _803 = _531 ? gnd : _802;
    assign _13 = _803;
    assign _492 = { _3891,
                    _13 };
    assign _832 = _221 ? _831 : gnd;
    assign _833 = _531 ? gnd : _832;
    assign _14 = _833;
    assign _489 = { _3891,
                    _14 };
    assign _862 = _221 ? _861 : gnd;
    assign _863 = _531 ? gnd : _862;
    assign _15 = _863;
    assign _486 = { _3891,
                    _15 };
    assign _892 = _221 ? _891 : gnd;
    assign _893 = _531 ? gnd : _892;
    assign _16 = _893;
    assign _483 = { _3891,
                    _16 };
    assign _922 = _221 ? _921 : gnd;
    assign _923 = _531 ? gnd : _922;
    assign _17 = _923;
    assign _480 = { _3891,
                    _17 };
    assign _952 = _221 ? _951 : gnd;
    assign _953 = _531 ? gnd : _952;
    assign _18 = _953;
    assign _477 = { _3891,
                    _18 };
    assign _982 = _221 ? _981 : gnd;
    assign _983 = _531 ? gnd : _982;
    assign _19 = _983;
    assign _474 = { _3891,
                    _19 };
    assign _1012 = _221 ? _1011 : gnd;
    assign _1013 = _531 ? gnd : _1012;
    assign _20 = _1013;
    assign _471 = { _3891,
                    _20 };
    assign _1031 = _221 ? _1030 : gnd;
    assign _1032 = _531 ? gnd : _1031;
    assign _21 = _1032;
    assign _468 = { _3891,
                    _21 };
    assign _1054 = _221 ? _1053 : gnd;
    assign _1055 = _531 ? gnd : _1054;
    assign _22 = _1055;
    assign _465 = { _3891,
                    _22 };
    assign _1084 = _221 ? _1083 : gnd;
    assign _1085 = _531 ? gnd : _1084;
    assign _23 = _1085;
    assign _462 = { _3891,
                    _23 };
    assign _1114 = _221 ? _1113 : gnd;
    assign _1115 = _531 ? gnd : _1114;
    assign _24 = _1115;
    assign _459 = { _3891,
                    _24 };
    assign _1144 = _221 ? _1143 : gnd;
    assign _1145 = _531 ? gnd : _1144;
    assign _25 = _1145;
    assign _456 = { _3891,
                    _25 };
    assign _1174 = _221 ? _1173 : gnd;
    assign _1175 = _531 ? gnd : _1174;
    assign _26 = _1175;
    assign _453 = { _3891,
                    _26 };
    assign _1204 = _221 ? _1203 : gnd;
    assign _1205 = _531 ? gnd : _1204;
    assign _27 = _1205;
    assign _450 = { _3891,
                    _27 };
    assign _1234 = _221 ? _1233 : gnd;
    assign _1235 = _531 ? gnd : _1234;
    assign _28 = _1235;
    assign _447 = { _3891,
                    _28 };
    assign _1264 = _221 ? _1263 : gnd;
    assign _1265 = _531 ? gnd : _1264;
    assign _29 = _1265;
    assign _444 = { _3891,
                    _29 };
    assign _1294 = _221 ? _1293 : gnd;
    assign _1295 = _531 ? gnd : _1294;
    assign _30 = _1295;
    assign _441 = { _3891,
                    _30 };
    assign _1313 = _221 ? _1312 : gnd;
    assign _1314 = _531 ? gnd : _1313;
    assign _31 = _1314;
    assign _438 = { _3891,
                    _31 };
    assign _1336 = _221 ? _1335 : gnd;
    assign _1337 = _531 ? gnd : _1336;
    assign _32 = _1337;
    assign _435 = { _3891,
                    _32 };
    assign _1366 = _221 ? _1365 : gnd;
    assign _1367 = _531 ? gnd : _1366;
    assign _33 = _1367;
    assign _432 = { _3891,
                    _33 };
    assign _1396 = _221 ? _1395 : gnd;
    assign _1397 = _531 ? gnd : _1396;
    assign _34 = _1397;
    assign _429 = { _3891,
                    _34 };
    assign _1426 = _221 ? _1425 : gnd;
    assign _1427 = _531 ? gnd : _1426;
    assign _35 = _1427;
    assign _426 = { _3891,
                    _35 };
    assign _1456 = _221 ? _1455 : gnd;
    assign _1457 = _531 ? gnd : _1456;
    assign _36 = _1457;
    assign _423 = { _3891,
                    _36 };
    assign _1486 = _221 ? _1485 : gnd;
    assign _1487 = _531 ? gnd : _1486;
    assign _37 = _1487;
    assign _420 = { _3891,
                    _37 };
    assign _1516 = _221 ? _1515 : gnd;
    assign _1517 = _531 ? gnd : _1516;
    assign _38 = _1517;
    assign _417 = { _3891,
                    _38 };
    assign _1546 = _221 ? _1545 : gnd;
    assign _1547 = _531 ? gnd : _1546;
    assign _39 = _1547;
    assign _414 = { _3891,
                    _39 };
    assign _1576 = _221 ? _1575 : gnd;
    assign _1577 = _531 ? gnd : _1576;
    assign _40 = _1577;
    assign _411 = { _3891,
                    _40 };
    assign _1595 = _221 ? _1594 : gnd;
    assign _1596 = _531 ? gnd : _1595;
    assign _41 = _1596;
    assign _408 = { _3891,
                    _41 };
    assign _1618 = _221 ? _1617 : gnd;
    assign _1619 = _531 ? gnd : _1618;
    assign _42 = _1619;
    assign _405 = { _3891,
                    _42 };
    assign _1648 = _221 ? _1647 : gnd;
    assign _1649 = _531 ? gnd : _1648;
    assign _43 = _1649;
    assign _402 = { _3891,
                    _43 };
    assign _1678 = _221 ? _1677 : gnd;
    assign _1679 = _531 ? gnd : _1678;
    assign _44 = _1679;
    assign _399 = { _3891,
                    _44 };
    assign _1708 = _221 ? _1707 : gnd;
    assign _1709 = _531 ? gnd : _1708;
    assign _45 = _1709;
    assign _396 = { _3891,
                    _45 };
    assign _1738 = _221 ? _1737 : gnd;
    assign _1739 = _531 ? gnd : _1738;
    assign _46 = _1739;
    assign _393 = { _3891,
                    _46 };
    assign _1768 = _221 ? _1767 : gnd;
    assign _1769 = _531 ? gnd : _1768;
    assign _47 = _1769;
    assign _390 = { _3891,
                    _47 };
    assign _1798 = _221 ? _1797 : gnd;
    assign _1799 = _531 ? gnd : _1798;
    assign _48 = _1799;
    assign _387 = { _3891,
                    _48 };
    assign _1828 = _221 ? _1827 : gnd;
    assign _1829 = _531 ? gnd : _1828;
    assign _49 = _1829;
    assign _384 = { _3891,
                    _49 };
    assign _1858 = _221 ? _1857 : gnd;
    assign _1859 = _531 ? gnd : _1858;
    assign _50 = _1859;
    assign _381 = { _3891,
                    _50 };
    assign _1877 = _221 ? _1876 : gnd;
    assign _1878 = _531 ? gnd : _1877;
    assign _51 = _1878;
    assign _378 = { _3891,
                    _51 };
    assign _1900 = _221 ? _1899 : gnd;
    assign _1901 = _531 ? gnd : _1900;
    assign _52 = _1901;
    assign _375 = { _3891,
                    _52 };
    assign _1930 = _221 ? _1929 : gnd;
    assign _1931 = _531 ? gnd : _1930;
    assign _53 = _1931;
    assign _372 = { _3891,
                    _53 };
    assign _1960 = _221 ? _1959 : gnd;
    assign _1961 = _531 ? gnd : _1960;
    assign _54 = _1961;
    assign _369 = { _3891,
                    _54 };
    assign _1990 = _221 ? _1989 : gnd;
    assign _1991 = _531 ? gnd : _1990;
    assign _55 = _1991;
    assign _366 = { _3891,
                    _55 };
    assign _2020 = _221 ? _2019 : gnd;
    assign _2021 = _531 ? gnd : _2020;
    assign _56 = _2021;
    assign _363 = { _3891,
                    _56 };
    assign _2050 = _221 ? _2049 : gnd;
    assign _2051 = _531 ? gnd : _2050;
    assign _57 = _2051;
    assign _360 = { _3891,
                    _57 };
    assign _2080 = _221 ? _2079 : gnd;
    assign _2081 = _531 ? gnd : _2080;
    assign _58 = _2081;
    assign _357 = { _3891,
                    _58 };
    assign _2110 = _221 ? _2109 : gnd;
    assign _2111 = _531 ? gnd : _2110;
    assign _59 = _2111;
    assign _354 = { _3891,
                    _59 };
    assign _2140 = _221 ? _2139 : gnd;
    assign _2141 = _531 ? gnd : _2140;
    assign _60 = _2141;
    assign _351 = { _3891,
                    _60 };
    assign _2159 = _221 ? _2158 : gnd;
    assign _2160 = _531 ? gnd : _2159;
    assign _61 = _2160;
    assign _348 = { _3891,
                    _61 };
    assign _2182 = _221 ? _2181 : gnd;
    assign _2183 = _531 ? gnd : _2182;
    assign _62 = _2183;
    assign _345 = { _3891,
                    _62 };
    assign _2212 = _221 ? _2211 : gnd;
    assign _2213 = _531 ? gnd : _2212;
    assign _63 = _2213;
    assign _342 = { _3891,
                    _63 };
    assign _2242 = _221 ? _2241 : gnd;
    assign _2243 = _531 ? gnd : _2242;
    assign _64 = _2243;
    assign _339 = { _3891,
                    _64 };
    assign _2272 = _221 ? _2271 : gnd;
    assign _2273 = _531 ? gnd : _2272;
    assign _65 = _2273;
    assign _336 = { _3891,
                    _65 };
    assign _2302 = _221 ? _2301 : gnd;
    assign _2303 = _531 ? gnd : _2302;
    assign _66 = _2303;
    assign _333 = { _3891,
                    _66 };
    assign _2332 = _221 ? _2331 : gnd;
    assign _2333 = _531 ? gnd : _2332;
    assign _67 = _2333;
    assign _330 = { _3891,
                    _67 };
    assign _2362 = _221 ? _2361 : gnd;
    assign _2363 = _531 ? gnd : _2362;
    assign _68 = _2363;
    assign _327 = { _3891,
                    _68 };
    assign _2392 = _221 ? _2391 : gnd;
    assign _2393 = _531 ? gnd : _2392;
    assign _69 = _2393;
    assign _324 = { _3891,
                    _69 };
    assign _2422 = _221 ? _2421 : gnd;
    assign _2423 = _531 ? gnd : _2422;
    assign _70 = _2423;
    assign _321 = { _3891,
                    _70 };
    assign _2441 = _221 ? _2440 : gnd;
    assign _2442 = _531 ? gnd : _2441;
    assign _71 = _2442;
    assign _318 = { _3891,
                    _71 };
    assign _2464 = _221 ? _2463 : gnd;
    assign _2465 = _531 ? gnd : _2464;
    assign _72 = _2465;
    assign _315 = { _3891,
                    _72 };
    assign _2494 = _221 ? _2493 : gnd;
    assign _2495 = _531 ? gnd : _2494;
    assign _73 = _2495;
    assign _312 = { _3891,
                    _73 };
    assign _2524 = _221 ? _2523 : gnd;
    assign _2525 = _531 ? gnd : _2524;
    assign _74 = _2525;
    assign _309 = { _3891,
                    _74 };
    assign _2554 = _221 ? _2553 : gnd;
    assign _2555 = _531 ? gnd : _2554;
    assign _75 = _2555;
    assign _306 = { _3891,
                    _75 };
    assign _2584 = _221 ? _2583 : gnd;
    assign _2585 = _531 ? gnd : _2584;
    assign _76 = _2585;
    assign _303 = { _3891,
                    _76 };
    assign _2614 = _221 ? _2613 : gnd;
    assign _2615 = _531 ? gnd : _2614;
    assign _77 = _2615;
    assign _300 = { _3891,
                    _77 };
    assign _2644 = _221 ? _2643 : gnd;
    assign _2645 = _531 ? gnd : _2644;
    assign _78 = _2645;
    assign _297 = { _3891,
                    _78 };
    assign _2674 = _221 ? _2673 : gnd;
    assign _2675 = _531 ? gnd : _2674;
    assign _79 = _2675;
    assign _294 = { _3891,
                    _79 };
    assign _2704 = _221 ? _2703 : gnd;
    assign _2705 = _531 ? gnd : _2704;
    assign _80 = _2705;
    assign _291 = { _3891,
                    _80 };
    assign _2723 = _221 ? _2722 : gnd;
    assign _2724 = _531 ? gnd : _2723;
    assign _81 = _2724;
    assign _288 = { _3891,
                    _81 };
    assign _2746 = _221 ? _2745 : gnd;
    assign _2747 = _531 ? gnd : _2746;
    assign _82 = _2747;
    assign _285 = { _3891,
                    _82 };
    assign _2776 = _221 ? _2775 : gnd;
    assign _2777 = _531 ? gnd : _2776;
    assign _83 = _2777;
    assign _282 = { _3891,
                    _83 };
    assign _2806 = _221 ? _2805 : gnd;
    assign _2807 = _531 ? gnd : _2806;
    assign _84 = _2807;
    assign _279 = { _3891,
                    _84 };
    assign _2836 = _221 ? _2835 : gnd;
    assign _2837 = _531 ? gnd : _2836;
    assign _85 = _2837;
    assign _276 = { _3891,
                    _85 };
    assign _2866 = _221 ? _2865 : gnd;
    assign _2867 = _531 ? gnd : _2866;
    assign _86 = _2867;
    assign _273 = { _3891,
                    _86 };
    assign _2896 = _221 ? _2895 : gnd;
    assign _2897 = _531 ? gnd : _2896;
    assign _87 = _2897;
    assign _270 = { _3891,
                    _87 };
    assign _2926 = _221 ? _2925 : gnd;
    assign _2927 = _531 ? gnd : _2926;
    assign _88 = _2927;
    assign _267 = { _3891,
                    _88 };
    assign _2956 = _221 ? _2955 : gnd;
    assign _2957 = _531 ? gnd : _2956;
    assign _89 = _2957;
    assign _264 = { _3891,
                    _89 };
    assign _2986 = _221 ? _2985 : gnd;
    assign _2987 = _531 ? gnd : _2986;
    assign _90 = _2987;
    assign _261 = { _3891,
                    _90 };
    assign _3005 = _221 ? _3004 : gnd;
    assign _3006 = _531 ? gnd : _3005;
    assign _91 = _3006;
    assign _258 = { _3891,
                    _91 };
    assign _3018 = _221 ? _3017 : gnd;
    assign _3019 = _531 ? gnd : _3018;
    assign _92 = _3019;
    assign _255 = { _3891,
                    _92 };
    assign _3037 = _221 ? _3036 : gnd;
    assign _3038 = _531 ? gnd : _3037;
    assign _93 = _3038;
    assign _252 = { _3891,
                    _93 };
    assign _3056 = _221 ? _3055 : gnd;
    assign _3057 = _531 ? gnd : _3056;
    assign _94 = _3057;
    assign _249 = { _3891,
                    _94 };
    assign _3075 = _221 ? _3074 : gnd;
    assign _3076 = _531 ? gnd : _3075;
    assign _95 = _3076;
    assign _246 = { _3891,
                    _95 };
    assign _3094 = _221 ? _3093 : gnd;
    assign _3095 = _531 ? gnd : _3094;
    assign _96 = _3095;
    assign _243 = { _3891,
                    _96 };
    assign _3113 = _221 ? _3112 : gnd;
    assign _3114 = _531 ? gnd : _3113;
    assign _97 = _3114;
    assign _240 = { _3891,
                    _97 };
    assign _3132 = _221 ? _3131 : gnd;
    assign _3133 = _531 ? gnd : _3132;
    assign _98 = _3133;
    assign _237 = { _3891,
                    _98 };
    assign _3151 = _221 ? _3150 : gnd;
    assign _3152 = _531 ? gnd : _3151;
    assign _99 = _3152;
    assign _234 = { _3891,
                    _99 };
    assign _3170 = _221 ? _3169 : gnd;
    assign _3171 = _531 ? gnd : _3170;
    assign _100 = _3171;
    assign _231 = { _3891,
                    _100 };
    assign _3576 = 4'b0100;
    assign _3573 = 3'b000;
    assign _3574 = { _3573,
                     _2648 };
    assign _3571 = { _3573,
                     _2678 };
    assign _2929 = 1'b0;
    assign _3165 = { _3573,
                     _2618 };
    assign _3162 = { _3573,
                     _2648 };
    assign _3159 = { _3573,
                     _2678 };
    assign _3146 = { _3573,
                     _2588 };
    assign _3143 = { _3573,
                     _2618 };
    assign _3140 = { _3573,
                     _2648 };
    assign _3127 = { _3573,
                     _2558 };
    assign _3124 = { _3573,
                     _2588 };
    assign _3121 = { _3573,
                     _2618 };
    assign _3108 = { _3573,
                     _2528 };
    assign _3105 = { _3573,
                     _2558 };
    assign _3102 = { _3573,
                     _2588 };
    assign _3089 = { _3573,
                     _2498 };
    assign _3086 = { _3573,
                     _2528 };
    assign _3083 = { _3573,
                     _2558 };
    assign _3070 = { _3573,
                     _2468 };
    assign _3067 = { _3573,
                     _2498 };
    assign _3064 = { _3573,
                     _2528 };
    assign _3051 = { _3573,
                     _2445 };
    assign _3048 = { _3573,
                     _2468 };
    assign _3045 = { _3573,
                     _2498 };
    assign _3032 = { _3573,
                     _2449 };
    assign _3029 = { _3573,
                     _2445 };
    assign _3026 = { _3573,
                     _2468 };
    assign _3013 = { _3573,
                     _2449 };
    assign _2771 = { _3573,
                     _2167 };
    assign _2768 = { _3573,
                     _2163 };
    assign _2765 = { _3573,
                     _2186 };
    assign _2762 = { _3573,
                     _2449 };
    assign _2801 = { _3573,
                     _2163 };
    assign _2798 = { _3573,
                     _2186 };
    assign _2795 = { _3573,
                     _2216 };
    assign _2792 = { _3573,
                     _2445 };
    assign _2831 = { _3573,
                     _2186 };
    assign _2828 = { _3573,
                     _2216 };
    assign _2825 = { _3573,
                     _2246 };
    assign _2822 = { _3573,
                     _2468 };
    assign _2861 = { _3573,
                     _2216 };
    assign _2858 = { _3573,
                     _2246 };
    assign _2855 = { _3573,
                     _2276 };
    assign _2852 = { _3573,
                     _2498 };
    assign _2891 = { _3573,
                     _2246 };
    assign _2888 = { _3573,
                     _2276 };
    assign _2885 = { _3573,
                     _2306 };
    assign _2882 = { _3573,
                     _2528 };
    assign _2921 = { _3573,
                     _2276 };
    assign _2918 = { _3573,
                     _2306 };
    assign _2915 = { _3573,
                     _2336 };
    assign _2912 = { _3573,
                     _2558 };
    assign _2951 = { _3573,
                     _2306 };
    assign _2948 = { _3573,
                     _2336 };
    assign _2945 = { _3573,
                     _2366 };
    assign _2942 = { _3573,
                     _2588 };
    assign _2981 = { _3573,
                     _2336 };
    assign _2978 = { _3573,
                     _2366 };
    assign _2975 = { _3573,
                     _2396 };
    assign _2972 = { _3573,
                     _2618 };
    assign _3000 = { _3573,
                     _2366 };
    assign _2718 = { _3573,
                     _2084 };
    assign _2715 = { _3573,
                     _2114 };
    assign _2699 = { _3573,
                     _2054 };
    assign _2696 = { _3573,
                     _2084 };
    assign _2693 = { _3573,
                     _2114 };
    assign _2669 = { _3573,
                     _2024 };
    assign _2666 = { _3573,
                     _2054 };
    assign _2663 = { _3573,
                     _2084 };
    assign _2639 = { _3573,
                     _1994 };
    assign _2636 = { _3573,
                     _2024 };
    assign _2633 = { _3573,
                     _2054 };
    assign _2609 = { _3573,
                     _1964 };
    assign _2606 = { _3573,
                     _1994 };
    assign _2603 = { _3573,
                     _2024 };
    assign _2579 = { _3573,
                     _1934 };
    assign _2576 = { _3573,
                     _1964 };
    assign _2573 = { _3573,
                     _1994 };
    assign _2549 = { _3573,
                     _1904 };
    assign _2546 = { _3573,
                     _1934 };
    assign _2543 = { _3573,
                     _1964 };
    assign _2519 = { _3573,
                     _1881 };
    assign _2516 = { _3573,
                     _1904 };
    assign _2513 = { _3573,
                     _1934 };
    assign _2489 = { _3573,
                     _1885 };
    assign _2486 = { _3573,
                     _1881 };
    assign _2483 = { _3573,
                     _1904 };
    assign _2480 = { _3573,
                     _2167 };
    assign _2477 = { _3573,
                     _2186 };
    assign _2459 = { _3573,
                     _1885 };
    assign _2207 = { _3573,
                     _1603 };
    assign _2204 = { _3573,
                     _1599 };
    assign _2201 = { _3573,
                     _1622 };
    assign _2198 = { _3573,
                     _1885 };
    assign _2237 = { _3573,
                     _1599 };
    assign _2234 = { _3573,
                     _1622 };
    assign _2231 = { _3573,
                     _1652 };
    assign _2228 = { _3573,
                     _1881 };
    assign _2267 = { _3573,
                     _1622 };
    assign _2264 = { _3573,
                     _1652 };
    assign _2261 = { _3573,
                     _1682 };
    assign _2258 = { _3573,
                     _1904 };
    assign _2297 = { _3573,
                     _1652 };
    assign _2294 = { _3573,
                     _1682 };
    assign _2291 = { _3573,
                     _1712 };
    assign _2288 = { _3573,
                     _1934 };
    assign _2327 = { _3573,
                     _1682 };
    assign _2324 = { _3573,
                     _1712 };
    assign _2321 = { _3573,
                     _1742 };
    assign _2318 = { _3573,
                     _1964 };
    assign _2357 = { _3573,
                     _1712 };
    assign _2354 = { _3573,
                     _1742 };
    assign _2351 = { _3573,
                     _1772 };
    assign _2348 = { _3573,
                     _1994 };
    assign _2387 = { _3573,
                     _1742 };
    assign _2384 = { _3573,
                     _1772 };
    assign _2381 = { _3573,
                     _1802 };
    assign _2378 = { _3573,
                     _2024 };
    assign _2417 = { _3573,
                     _1772 };
    assign _2414 = { _3573,
                     _1802 };
    assign _2411 = { _3573,
                     _1832 };
    assign _2408 = { _3573,
                     _2054 };
    assign _2436 = { _3573,
                     _1802 };
    assign _2154 = { _3573,
                     _1520 };
    assign _2151 = { _3573,
                     _1550 };
    assign _2135 = { _3573,
                     _1490 };
    assign _2132 = { _3573,
                     _1520 };
    assign _2129 = { _3573,
                     _1550 };
    assign _2105 = { _3573,
                     _1460 };
    assign _2102 = { _3573,
                     _1490 };
    assign _2099 = { _3573,
                     _1520 };
    assign _2075 = { _3573,
                     _1430 };
    assign _2072 = { _3573,
                     _1460 };
    assign _2069 = { _3573,
                     _1490 };
    assign _2045 = { _3573,
                     _1400 };
    assign _2042 = { _3573,
                     _1430 };
    assign _2039 = { _3573,
                     _1460 };
    assign _2015 = { _3573,
                     _1370 };
    assign _2012 = { _3573,
                     _1400 };
    assign _2009 = { _3573,
                     _1430 };
    assign _1985 = { _3573,
                     _1340 };
    assign _1982 = { _3573,
                     _1370 };
    assign _1979 = { _3573,
                     _1400 };
    assign _1955 = { _3573,
                     _1317 };
    assign _1952 = { _3573,
                     _1340 };
    assign _1949 = { _3573,
                     _1370 };
    assign _1925 = { _3573,
                     _1321 };
    assign _1922 = { _3573,
                     _1317 };
    assign _1919 = { _3573,
                     _1340 };
    assign _1916 = { _3573,
                     _1603 };
    assign _1913 = { _3573,
                     _1622 };
    assign _1895 = { _3573,
                     _1321 };
    assign _1643 = { _3573,
                     _1039 };
    assign _1640 = { _3573,
                     _1035 };
    assign _1637 = { _3573,
                     _1058 };
    assign _1634 = { _3573,
                     _1321 };
    assign _1673 = { _3573,
                     _1035 };
    assign _1670 = { _3573,
                     _1058 };
    assign _1667 = { _3573,
                     _1088 };
    assign _1664 = { _3573,
                     _1317 };
    assign _1703 = { _3573,
                     _1058 };
    assign _1700 = { _3573,
                     _1088 };
    assign _1697 = { _3573,
                     _1118 };
    assign _1694 = { _3573,
                     _1340 };
    assign _1733 = { _3573,
                     _1088 };
    assign _1730 = { _3573,
                     _1118 };
    assign _1727 = { _3573,
                     _1148 };
    assign _1724 = { _3573,
                     _1370 };
    assign _1763 = { _3573,
                     _1118 };
    assign _1760 = { _3573,
                     _1148 };
    assign _1757 = { _3573,
                     _1178 };
    assign _1754 = { _3573,
                     _1400 };
    assign _1793 = { _3573,
                     _1148 };
    assign _1790 = { _3573,
                     _1178 };
    assign _1787 = { _3573,
                     _1208 };
    assign _1784 = { _3573,
                     _1430 };
    assign _1823 = { _3573,
                     _1178 };
    assign _1820 = { _3573,
                     _1208 };
    assign _1817 = { _3573,
                     _1238 };
    assign _1814 = { _3573,
                     _1460 };
    assign _1853 = { _3573,
                     _1208 };
    assign _1850 = { _3573,
                     _1238 };
    assign _1847 = { _3573,
                     _1268 };
    assign _1844 = { _3573,
                     _1490 };
    assign _1872 = { _3573,
                     _1238 };
    assign _1590 = { _3573,
                     _956 };
    assign _1587 = { _3573,
                     _986 };
    assign _1571 = { _3573,
                     _926 };
    assign _1568 = { _3573,
                     _956 };
    assign _1565 = { _3573,
                     _986 };
    assign _1541 = { _3573,
                     _896 };
    assign _1538 = { _3573,
                     _926 };
    assign _1535 = { _3573,
                     _956 };
    assign _1511 = { _3573,
                     _866 };
    assign _1508 = { _3573,
                     _896 };
    assign _1505 = { _3573,
                     _926 };
    assign _1481 = { _3573,
                     _836 };
    assign _1478 = { _3573,
                     _866 };
    assign _1475 = { _3573,
                     _896 };
    assign _1451 = { _3573,
                     _806 };
    assign _1448 = { _3573,
                     _836 };
    assign _1445 = { _3573,
                     _866 };
    assign _1421 = { _3573,
                     _776 };
    assign _1418 = { _3573,
                     _806 };
    assign _1415 = { _3573,
                     _836 };
    assign _1391 = { _3573,
                     _753 };
    assign _1388 = { _3573,
                     _776 };
    assign _1385 = { _3573,
                     _806 };
    assign _1361 = { _3573,
                     _757 };
    assign _1358 = { _3573,
                     _753 };
    assign _1355 = { _3573,
                     _776 };
    assign _1352 = { _3573,
                     _1039 };
    assign _1349 = { _3573,
                     _1058 };
    assign _1331 = { _3573,
                     _757 };
    assign _1079 = { _3573,
                     _541 };
    assign _1076 = { _3573,
                     _537 };
    assign _1073 = { _3573,
                     _556 };
    assign _1070 = { _3573,
                     _757 };
    assign _1109 = { _3573,
                     _537 };
    assign _1106 = { _3573,
                     _556 };
    assign _1103 = { _3573,
                     _579 };
    assign _1100 = { _3573,
                     _753 };
    assign _1139 = { _3573,
                     _556 };
    assign _1136 = { _3573,
                     _579 };
    assign _1133 = { _3573,
                     _602 };
    assign _1130 = { _3573,
                     _776 };
    assign _1169 = { _3573,
                     _579 };
    assign _1166 = { _3573,
                     _602 };
    assign _1163 = { _3573,
                     _625 };
    assign _1160 = { _3573,
                     _806 };
    assign _1199 = { _3573,
                     _602 };
    assign _1196 = { _3573,
                     _625 };
    assign _1193 = { _3573,
                     _648 };
    assign _1190 = { _3573,
                     _836 };
    assign _1229 = { _3573,
                     _625 };
    assign _1226 = { _3573,
                     _648 };
    assign _1223 = { _3573,
                     _671 };
    assign _1220 = { _3573,
                     _866 };
    assign _1259 = { _3573,
                     _648 };
    assign _1256 = { _3573,
                     _671 };
    assign _1253 = { _3573,
                     _694 };
    assign _1250 = { _3573,
                     _896 };
    assign _1289 = { _3573,
                     _671 };
    assign _1286 = { _3573,
                     _694 };
    assign _1283 = { _3573,
                     _717 };
    assign _1280 = { _3573,
                     _926 };
    assign _1308 = { _3573,
                     _694 };
    assign _1026 = { _3573,
                     _704 };
    assign _1023 = { _3573,
                     _727 };
    assign _1007 = { _3573,
                     _681 };
    assign _1004 = { _3573,
                     _704 };
    assign _1001 = { _3573,
                     _727 };
    assign _977 = { _3573,
                    _658 };
    assign _974 = { _3573,
                    _681 };
    assign _971 = { _3573,
                    _704 };
    assign _947 = { _3573,
                    _635 };
    assign _944 = { _3573,
                    _658 };
    assign _941 = { _3573,
                    _681 };
    assign _917 = { _3573,
                    _612 };
    assign _914 = { _3573,
                    _635 };
    assign _911 = { _3573,
                    _658 };
    assign _887 = { _3573,
                    _589 };
    assign _884 = { _3573,
                    _612 };
    assign _881 = { _3573,
                    _635 };
    assign _857 = { _3573,
                    _566 };
    assign _854 = { _3573,
                    _589 };
    assign _851 = { _3573,
                    _612 };
    assign _827 = { _3573,
                    _546 };
    assign _824 = { _3573,
                    _566 };
    assign _821 = { _3573,
                    _589 };
    assign _797 = { _3573,
                    _534 };
    assign _794 = { _3573,
                    _546 };
    assign _791 = { _3573,
                    _566 };
    assign _788 = { _3573,
                    _541 };
    assign _785 = { _3573,
                    _556 };
    assign _767 = { _3573,
                    _534 };
    assign _547 = { _3573,
                    _546 };
    assign _542 = { _3573,
                    _541 };
    assign _538 = { _3573,
                    _537 };
    assign _543 = _538 + _542;
    assign _548 = _543 + _547;
    assign _550 = _548 < _3576;
    assign _551 = _534 & _550;
    assign _3172 = ~ _551;
    assign _3173 = _534 & _3172;
    assign _3174 = _221 ? _3173 : _534;
    assign _3175 = _531 ? _546 : _3174;
    assign _101 = _3175;
    always @(posedge _209) begin
        if (_223)
            _534 <= _2929;
        else
            _534 <= _101;
    end
    assign _570 = { _3573,
                    _534 };
    assign _593 = { _3573,
                    _546 };
    assign _616 = { _3573,
                    _566 };
    assign _639 = { _3573,
                    _589 };
    assign _662 = { _3573,
                    _612 };
    assign _685 = { _3573,
                    _635 };
    assign _708 = { _3573,
                    _658 };
    assign _731 = { _3573,
                    _681 };
    assign _744 = { _3573,
                    _704 };
    assign _741 = { _3573,
                    _694 };
    assign _739 = { _3573,
                    _717 };
    assign _742 = _739 + _741;
    assign _745 = _742 + _744;
    assign _747 = _745 < _3576;
    assign _748 = _727 & _747;
    assign _3176 = ~ _748;
    assign _3177 = _727 & _3176;
    assign _3178 = _221 ? _3177 : _727;
    assign _3179 = _531 ? _541 : _3178;
    assign _102 = _3179;
    always @(posedge _209) begin
        if (_223)
            _727 <= _2929;
        else
            _727 <= _102;
    end
    assign _728 = { _3573,
                    _727 };
    assign _723 = { _3573,
                    _671 };
    assign _720 = { _3573,
                    _694 };
    assign _718 = { _3573,
                    _717 };
    assign _721 = _718 + _720;
    assign _724 = _721 + _723;
    assign _729 = _724 + _728;
    assign _732 = _729 + _731;
    assign _734 = _732 < _3576;
    assign _735 = _704 & _734;
    assign _3180 = ~ _735;
    assign _3181 = _704 & _3180;
    assign _3182 = _221 ? _3181 : _704;
    assign _3183 = _531 ? _727 : _3182;
    assign _103 = _3183;
    always @(posedge _209) begin
        if (_223)
            _704 <= _2929;
        else
            _704 <= _103;
    end
    assign _705 = { _3573,
                    _704 };
    assign _700 = { _3573,
                    _648 };
    assign _697 = { _3573,
                    _671 };
    assign _695 = { _3573,
                    _694 };
    assign _698 = _695 + _697;
    assign _701 = _698 + _700;
    assign _706 = _701 + _705;
    assign _709 = _706 + _708;
    assign _711 = _709 < _3576;
    assign _712 = _681 & _711;
    assign _3184 = ~ _712;
    assign _3185 = _681 & _3184;
    assign _3186 = _221 ? _3185 : _681;
    assign _3187 = _531 ? _704 : _3186;
    assign _104 = _3187;
    always @(posedge _209) begin
        if (_223)
            _681 <= _2929;
        else
            _681 <= _104;
    end
    assign _682 = { _3573,
                    _681 };
    assign _677 = { _3573,
                    _625 };
    assign _674 = { _3573,
                    _648 };
    assign _672 = { _3573,
                    _671 };
    assign _675 = _672 + _674;
    assign _678 = _675 + _677;
    assign _683 = _678 + _682;
    assign _686 = _683 + _685;
    assign _688 = _686 < _3576;
    assign _689 = _658 & _688;
    assign _3188 = ~ _689;
    assign _3189 = _658 & _3188;
    assign _3190 = _221 ? _3189 : _658;
    assign _3191 = _531 ? _681 : _3190;
    assign _105 = _3191;
    always @(posedge _209) begin
        if (_223)
            _658 <= _2929;
        else
            _658 <= _105;
    end
    assign _659 = { _3573,
                    _658 };
    assign _654 = { _3573,
                    _602 };
    assign _651 = { _3573,
                    _625 };
    assign _649 = { _3573,
                    _648 };
    assign _652 = _649 + _651;
    assign _655 = _652 + _654;
    assign _660 = _655 + _659;
    assign _663 = _660 + _662;
    assign _665 = _663 < _3576;
    assign _666 = _635 & _665;
    assign _3192 = ~ _666;
    assign _3193 = _635 & _3192;
    assign _3194 = _221 ? _3193 : _635;
    assign _3195 = _531 ? _658 : _3194;
    assign _106 = _3195;
    always @(posedge _209) begin
        if (_223)
            _635 <= _2929;
        else
            _635 <= _106;
    end
    assign _636 = { _3573,
                    _635 };
    assign _631 = { _3573,
                    _579 };
    assign _628 = { _3573,
                    _602 };
    assign _626 = { _3573,
                    _625 };
    assign _629 = _626 + _628;
    assign _632 = _629 + _631;
    assign _637 = _632 + _636;
    assign _640 = _637 + _639;
    assign _642 = _640 < _3576;
    assign _643 = _612 & _642;
    assign _3196 = ~ _643;
    assign _3197 = _612 & _3196;
    assign _3198 = _221 ? _3197 : _612;
    assign _3199 = _531 ? _635 : _3198;
    assign _107 = _3199;
    always @(posedge _209) begin
        if (_223)
            _612 <= _2929;
        else
            _612 <= _107;
    end
    assign _613 = { _3573,
                    _612 };
    assign _608 = { _3573,
                    _556 };
    assign _605 = { _3573,
                    _579 };
    assign _603 = { _3573,
                    _602 };
    assign _606 = _603 + _605;
    assign _609 = _606 + _608;
    assign _614 = _609 + _613;
    assign _617 = _614 + _616;
    assign _619 = _617 < _3576;
    assign _620 = _589 & _619;
    assign _3200 = ~ _620;
    assign _3201 = _589 & _3200;
    assign _3202 = _221 ? _3201 : _589;
    assign _3203 = _531 ? _612 : _3202;
    assign _108 = _3203;
    always @(posedge _209) begin
        if (_223)
            _589 <= _2929;
        else
            _589 <= _108;
    end
    assign _590 = { _3573,
                    _589 };
    assign _585 = { _3573,
                    _537 };
    assign _582 = { _3573,
                    _556 };
    assign _580 = { _3573,
                    _579 };
    assign _583 = _580 + _582;
    assign _586 = _583 + _585;
    assign _591 = _586 + _590;
    assign _594 = _591 + _593;
    assign _596 = _594 < _3576;
    assign _597 = _566 & _596;
    assign _3204 = ~ _597;
    assign _3205 = _566 & _3204;
    assign _3206 = _221 ? _3205 : _566;
    assign _3207 = _531 ? _589 : _3206;
    assign _109 = _3207;
    always @(posedge _209) begin
        if (_223)
            _566 <= _2929;
        else
            _566 <= _109;
    end
    assign _567 = { _3573,
                    _566 };
    assign _562 = { _3573,
                    _541 };
    assign _559 = { _3573,
                    _537 };
    assign _557 = { _3573,
                    _556 };
    assign _560 = _557 + _559;
    assign _563 = _560 + _562;
    assign _568 = _563 + _567;
    assign _571 = _568 + _570;
    assign _573 = _571 < _3576;
    assign _574 = _546 & _573;
    assign _3208 = ~ _574;
    assign _3209 = _546 & _3208;
    assign _3210 = _221 ? _3209 : _546;
    assign _3211 = _531 ? _566 : _3210;
    assign _110 = _3211;
    always @(posedge _209) begin
        if (_223)
            _546 <= _2929;
        else
            _546 <= _110;
    end
    assign _764 = { _3573,
                    _546 };
    assign _761 = { _3573,
                    _537 };
    assign _758 = { _3573,
                    _757 };
    assign _754 = { _3573,
                    _753 };
    assign _759 = _754 + _758;
    assign _762 = _759 + _761;
    assign _765 = _762 + _764;
    assign _768 = _765 + _767;
    assign _770 = _768 < _3576;
    assign _771 = _541 & _770;
    assign _3212 = ~ _771;
    assign _3213 = _541 & _3212;
    assign _3214 = _221 ? _3213 : _541;
    assign _3215 = _531 ? _537 : _3214;
    assign _111 = _3215;
    always @(posedge _209) begin
        if (_223)
            _541 <= _2929;
        else
            _541 <= _111;
    end
    assign _1049 = { _3573,
                     _541 };
    assign _1046 = { _3573,
                     _537 };
    assign _1043 = { _3573,
                     _753 };
    assign _1040 = { _3573,
                     _1039 };
    assign _1036 = { _3573,
                     _1035 };
    assign _1041 = _1036 + _1040;
    assign _1044 = _1041 + _1043;
    assign _1047 = _1044 + _1046;
    assign _1050 = _1047 + _1049;
    assign _1052 = _1050 < _3576;
    assign _1053 = _757 & _1052;
    assign _3216 = ~ _1053;
    assign _3217 = _757 & _3216;
    assign _3218 = _221 ? _3217 : _757;
    assign _3219 = _531 ? _753 : _3218;
    assign _112 = _3219;
    always @(posedge _209) begin
        if (_223)
            _757 <= _2929;
        else
            _757 <= _112;
    end
    assign _782 = { _3573,
                    _757 };
    assign _779 = { _3573,
                    _753 };
    assign _777 = { _3573,
                    _776 };
    assign _780 = _777 + _779;
    assign _783 = _780 + _782;
    assign _786 = _783 + _785;
    assign _789 = _786 + _788;
    assign _792 = _789 + _791;
    assign _795 = _792 + _794;
    assign _798 = _795 + _797;
    assign _800 = _798 < _3576;
    assign _801 = _537 & _800;
    assign _3220 = ~ _801;
    assign _3221 = _537 & _3220;
    assign _3222 = _221 ? _3221 : _537;
    assign _3223 = _531 ? _556 : _3222;
    assign _113 = _3223;
    always @(posedge _209) begin
        if (_223)
            _537 <= _2929;
        else
            _537 <= _113;
    end
    assign _818 = { _3573,
                    _537 };
    assign _815 = { _3573,
                    _579 };
    assign _812 = { _3573,
                    _753 };
    assign _809 = { _3573,
                    _776 };
    assign _807 = { _3573,
                    _806 };
    assign _810 = _807 + _809;
    assign _813 = _810 + _812;
    assign _816 = _813 + _815;
    assign _819 = _816 + _818;
    assign _822 = _819 + _821;
    assign _825 = _822 + _824;
    assign _828 = _825 + _827;
    assign _830 = _828 < _3576;
    assign _831 = _556 & _830;
    assign _3224 = ~ _831;
    assign _3225 = _556 & _3224;
    assign _3226 = _221 ? _3225 : _556;
    assign _3227 = _531 ? _579 : _3226;
    assign _114 = _3227;
    always @(posedge _209) begin
        if (_223)
            _556 <= _2929;
        else
            _556 <= _114;
    end
    assign _848 = { _3573,
                    _556 };
    assign _845 = { _3573,
                    _602 };
    assign _842 = { _3573,
                    _776 };
    assign _839 = { _3573,
                    _806 };
    assign _837 = { _3573,
                    _836 };
    assign _840 = _837 + _839;
    assign _843 = _840 + _842;
    assign _846 = _843 + _845;
    assign _849 = _846 + _848;
    assign _852 = _849 + _851;
    assign _855 = _852 + _854;
    assign _858 = _855 + _857;
    assign _860 = _858 < _3576;
    assign _861 = _579 & _860;
    assign _3228 = ~ _861;
    assign _3229 = _579 & _3228;
    assign _3230 = _221 ? _3229 : _579;
    assign _3231 = _531 ? _602 : _3230;
    assign _115 = _3231;
    always @(posedge _209) begin
        if (_223)
            _579 <= _2929;
        else
            _579 <= _115;
    end
    assign _878 = { _3573,
                    _579 };
    assign _875 = { _3573,
                    _625 };
    assign _872 = { _3573,
                    _806 };
    assign _869 = { _3573,
                    _836 };
    assign _867 = { _3573,
                    _866 };
    assign _870 = _867 + _869;
    assign _873 = _870 + _872;
    assign _876 = _873 + _875;
    assign _879 = _876 + _878;
    assign _882 = _879 + _881;
    assign _885 = _882 + _884;
    assign _888 = _885 + _887;
    assign _890 = _888 < _3576;
    assign _891 = _602 & _890;
    assign _3232 = ~ _891;
    assign _3233 = _602 & _3232;
    assign _3234 = _221 ? _3233 : _602;
    assign _3235 = _531 ? _625 : _3234;
    assign _116 = _3235;
    always @(posedge _209) begin
        if (_223)
            _602 <= _2929;
        else
            _602 <= _116;
    end
    assign _908 = { _3573,
                    _602 };
    assign _905 = { _3573,
                    _648 };
    assign _902 = { _3573,
                    _836 };
    assign _899 = { _3573,
                    _866 };
    assign _897 = { _3573,
                    _896 };
    assign _900 = _897 + _899;
    assign _903 = _900 + _902;
    assign _906 = _903 + _905;
    assign _909 = _906 + _908;
    assign _912 = _909 + _911;
    assign _915 = _912 + _914;
    assign _918 = _915 + _917;
    assign _920 = _918 < _3576;
    assign _921 = _625 & _920;
    assign _3236 = ~ _921;
    assign _3237 = _625 & _3236;
    assign _3238 = _221 ? _3237 : _625;
    assign _3239 = _531 ? _648 : _3238;
    assign _117 = _3239;
    always @(posedge _209) begin
        if (_223)
            _625 <= _2929;
        else
            _625 <= _117;
    end
    assign _938 = { _3573,
                    _625 };
    assign _935 = { _3573,
                    _671 };
    assign _932 = { _3573,
                    _866 };
    assign _929 = { _3573,
                    _896 };
    assign _927 = { _3573,
                    _926 };
    assign _930 = _927 + _929;
    assign _933 = _930 + _932;
    assign _936 = _933 + _935;
    assign _939 = _936 + _938;
    assign _942 = _939 + _941;
    assign _945 = _942 + _944;
    assign _948 = _945 + _947;
    assign _950 = _948 < _3576;
    assign _951 = _648 & _950;
    assign _3240 = ~ _951;
    assign _3241 = _648 & _3240;
    assign _3242 = _221 ? _3241 : _648;
    assign _3243 = _531 ? _671 : _3242;
    assign _118 = _3243;
    always @(posedge _209) begin
        if (_223)
            _648 <= _2929;
        else
            _648 <= _118;
    end
    assign _968 = { _3573,
                    _648 };
    assign _965 = { _3573,
                    _694 };
    assign _962 = { _3573,
                    _896 };
    assign _959 = { _3573,
                    _926 };
    assign _957 = { _3573,
                    _956 };
    assign _960 = _957 + _959;
    assign _963 = _960 + _962;
    assign _966 = _963 + _965;
    assign _969 = _966 + _968;
    assign _972 = _969 + _971;
    assign _975 = _972 + _974;
    assign _978 = _975 + _977;
    assign _980 = _978 < _3576;
    assign _981 = _671 & _980;
    assign _3244 = ~ _981;
    assign _3245 = _671 & _3244;
    assign _3246 = _221 ? _3245 : _671;
    assign _3247 = _531 ? _694 : _3246;
    assign _119 = _3247;
    always @(posedge _209) begin
        if (_223)
            _671 <= _2929;
        else
            _671 <= _119;
    end
    assign _998 = { _3573,
                    _671 };
    assign _995 = { _3573,
                    _717 };
    assign _992 = { _3573,
                    _926 };
    assign _989 = { _3573,
                    _956 };
    assign _987 = { _3573,
                    _986 };
    assign _990 = _987 + _989;
    assign _993 = _990 + _992;
    assign _996 = _993 + _995;
    assign _999 = _996 + _998;
    assign _1002 = _999 + _1001;
    assign _1005 = _1002 + _1004;
    assign _1008 = _1005 + _1007;
    assign _1010 = _1008 < _3576;
    assign _1011 = _694 & _1010;
    assign _3248 = ~ _1011;
    assign _3249 = _694 & _3248;
    assign _3250 = _221 ? _3249 : _694;
    assign _3251 = _531 ? _717 : _3250;
    assign _120 = _3251;
    always @(posedge _209) begin
        if (_223)
            _694 <= _2929;
        else
            _694 <= _120;
    end
    assign _1020 = { _3573,
                     _694 };
    assign _1017 = { _3573,
                     _956 };
    assign _1015 = { _3573,
                     _986 };
    assign _1018 = _1015 + _1017;
    assign _1021 = _1018 + _1020;
    assign _1024 = _1021 + _1023;
    assign _1027 = _1024 + _1026;
    assign _1029 = _1027 < _3576;
    assign _1030 = _717 & _1029;
    assign _3252 = ~ _1030;
    assign _3253 = _717 & _3252;
    assign _3254 = _221 ? _3253 : _717;
    assign _3255 = _531 ? _757 : _3254;
    assign _121 = _3255;
    always @(posedge _209) begin
        if (_223)
            _717 <= _2929;
        else
            _717 <= _121;
    end
    assign _1305 = { _3573,
                     _717 };
    assign _1302 = { _3573,
                     _956 };
    assign _1299 = { _3573,
                     _1238 };
    assign _1297 = { _3573,
                     _1268 };
    assign _1300 = _1297 + _1299;
    assign _1303 = _1300 + _1302;
    assign _1306 = _1303 + _1305;
    assign _1309 = _1306 + _1308;
    assign _1311 = _1309 < _3576;
    assign _1312 = _986 & _1311;
    assign _3256 = ~ _1312;
    assign _3257 = _986 & _3256;
    assign _3258 = _221 ? _3257 : _986;
    assign _3259 = _531 ? _1039 : _3258;
    assign _122 = _3259;
    always @(posedge _209) begin
        if (_223)
            _986 <= _2929;
        else
            _986 <= _122;
    end
    assign _1277 = { _3573,
                     _986 };
    assign _1274 = { _3573,
                     _1208 };
    assign _1271 = { _3573,
                     _1238 };
    assign _1269 = { _3573,
                     _1268 };
    assign _1272 = _1269 + _1271;
    assign _1275 = _1272 + _1274;
    assign _1278 = _1275 + _1277;
    assign _1281 = _1278 + _1280;
    assign _1284 = _1281 + _1283;
    assign _1287 = _1284 + _1286;
    assign _1290 = _1287 + _1289;
    assign _1292 = _1290 < _3576;
    assign _1293 = _956 & _1292;
    assign _3260 = ~ _1293;
    assign _3261 = _956 & _3260;
    assign _3262 = _221 ? _3261 : _956;
    assign _3263 = _531 ? _986 : _3262;
    assign _123 = _3263;
    always @(posedge _209) begin
        if (_223)
            _956 <= _2929;
        else
            _956 <= _123;
    end
    assign _1247 = { _3573,
                     _956 };
    assign _1244 = { _3573,
                     _1178 };
    assign _1241 = { _3573,
                     _1208 };
    assign _1239 = { _3573,
                     _1238 };
    assign _1242 = _1239 + _1241;
    assign _1245 = _1242 + _1244;
    assign _1248 = _1245 + _1247;
    assign _1251 = _1248 + _1250;
    assign _1254 = _1251 + _1253;
    assign _1257 = _1254 + _1256;
    assign _1260 = _1257 + _1259;
    assign _1262 = _1260 < _3576;
    assign _1263 = _926 & _1262;
    assign _3264 = ~ _1263;
    assign _3265 = _926 & _3264;
    assign _3266 = _221 ? _3265 : _926;
    assign _3267 = _531 ? _956 : _3266;
    assign _124 = _3267;
    always @(posedge _209) begin
        if (_223)
            _926 <= _2929;
        else
            _926 <= _124;
    end
    assign _1217 = { _3573,
                     _926 };
    assign _1214 = { _3573,
                     _1148 };
    assign _1211 = { _3573,
                     _1178 };
    assign _1209 = { _3573,
                     _1208 };
    assign _1212 = _1209 + _1211;
    assign _1215 = _1212 + _1214;
    assign _1218 = _1215 + _1217;
    assign _1221 = _1218 + _1220;
    assign _1224 = _1221 + _1223;
    assign _1227 = _1224 + _1226;
    assign _1230 = _1227 + _1229;
    assign _1232 = _1230 < _3576;
    assign _1233 = _896 & _1232;
    assign _3268 = ~ _1233;
    assign _3269 = _896 & _3268;
    assign _3270 = _221 ? _3269 : _896;
    assign _3271 = _531 ? _926 : _3270;
    assign _125 = _3271;
    always @(posedge _209) begin
        if (_223)
            _896 <= _2929;
        else
            _896 <= _125;
    end
    assign _1187 = { _3573,
                     _896 };
    assign _1184 = { _3573,
                     _1118 };
    assign _1181 = { _3573,
                     _1148 };
    assign _1179 = { _3573,
                     _1178 };
    assign _1182 = _1179 + _1181;
    assign _1185 = _1182 + _1184;
    assign _1188 = _1185 + _1187;
    assign _1191 = _1188 + _1190;
    assign _1194 = _1191 + _1193;
    assign _1197 = _1194 + _1196;
    assign _1200 = _1197 + _1199;
    assign _1202 = _1200 < _3576;
    assign _1203 = _866 & _1202;
    assign _3272 = ~ _1203;
    assign _3273 = _866 & _3272;
    assign _3274 = _221 ? _3273 : _866;
    assign _3275 = _531 ? _896 : _3274;
    assign _126 = _3275;
    always @(posedge _209) begin
        if (_223)
            _866 <= _2929;
        else
            _866 <= _126;
    end
    assign _1157 = { _3573,
                     _866 };
    assign _1154 = { _3573,
                     _1088 };
    assign _1151 = { _3573,
                     _1118 };
    assign _1149 = { _3573,
                     _1148 };
    assign _1152 = _1149 + _1151;
    assign _1155 = _1152 + _1154;
    assign _1158 = _1155 + _1157;
    assign _1161 = _1158 + _1160;
    assign _1164 = _1161 + _1163;
    assign _1167 = _1164 + _1166;
    assign _1170 = _1167 + _1169;
    assign _1172 = _1170 < _3576;
    assign _1173 = _836 & _1172;
    assign _3276 = ~ _1173;
    assign _3277 = _836 & _3276;
    assign _3278 = _221 ? _3277 : _836;
    assign _3279 = _531 ? _866 : _3278;
    assign _127 = _3279;
    always @(posedge _209) begin
        if (_223)
            _836 <= _2929;
        else
            _836 <= _127;
    end
    assign _1127 = { _3573,
                     _836 };
    assign _1124 = { _3573,
                     _1058 };
    assign _1121 = { _3573,
                     _1088 };
    assign _1119 = { _3573,
                     _1118 };
    assign _1122 = _1119 + _1121;
    assign _1125 = _1122 + _1124;
    assign _1128 = _1125 + _1127;
    assign _1131 = _1128 + _1130;
    assign _1134 = _1131 + _1133;
    assign _1137 = _1134 + _1136;
    assign _1140 = _1137 + _1139;
    assign _1142 = _1140 < _3576;
    assign _1143 = _806 & _1142;
    assign _3280 = ~ _1143;
    assign _3281 = _806 & _3280;
    assign _3282 = _221 ? _3281 : _806;
    assign _3283 = _531 ? _836 : _3282;
    assign _128 = _3283;
    always @(posedge _209) begin
        if (_223)
            _806 <= _2929;
        else
            _806 <= _128;
    end
    assign _1097 = { _3573,
                     _806 };
    assign _1094 = { _3573,
                     _1035 };
    assign _1091 = { _3573,
                     _1058 };
    assign _1089 = { _3573,
                     _1088 };
    assign _1092 = _1089 + _1091;
    assign _1095 = _1092 + _1094;
    assign _1098 = _1095 + _1097;
    assign _1101 = _1098 + _1100;
    assign _1104 = _1101 + _1103;
    assign _1107 = _1104 + _1106;
    assign _1110 = _1107 + _1109;
    assign _1112 = _1110 < _3576;
    assign _1113 = _776 & _1112;
    assign _3284 = ~ _1113;
    assign _3285 = _776 & _3284;
    assign _3286 = _221 ? _3285 : _776;
    assign _3287 = _531 ? _806 : _3286;
    assign _129 = _3287;
    always @(posedge _209) begin
        if (_223)
            _776 <= _2929;
        else
            _776 <= _129;
    end
    assign _1067 = { _3573,
                     _776 };
    assign _1064 = { _3573,
                     _1039 };
    assign _1061 = { _3573,
                     _1035 };
    assign _1059 = { _3573,
                     _1058 };
    assign _1062 = _1059 + _1061;
    assign _1065 = _1062 + _1064;
    assign _1068 = _1065 + _1067;
    assign _1071 = _1068 + _1070;
    assign _1074 = _1071 + _1073;
    assign _1077 = _1074 + _1076;
    assign _1080 = _1077 + _1079;
    assign _1082 = _1080 < _3576;
    assign _1083 = _753 & _1082;
    assign _3288 = ~ _1083;
    assign _3289 = _753 & _3288;
    assign _3290 = _221 ? _3289 : _753;
    assign _3291 = _531 ? _776 : _3290;
    assign _130 = _3291;
    always @(posedge _209) begin
        if (_223)
            _753 <= _2929;
        else
            _753 <= _130;
    end
    assign _1328 = { _3573,
                     _753 };
    assign _1325 = { _3573,
                     _1035 };
    assign _1322 = { _3573,
                     _1321 };
    assign _1318 = { _3573,
                     _1317 };
    assign _1323 = _1318 + _1322;
    assign _1326 = _1323 + _1325;
    assign _1329 = _1326 + _1328;
    assign _1332 = _1329 + _1331;
    assign _1334 = _1332 < _3576;
    assign _1335 = _1039 & _1334;
    assign _3292 = ~ _1335;
    assign _3293 = _1039 & _3292;
    assign _3294 = _221 ? _3293 : _1039;
    assign _3295 = _531 ? _1035 : _3294;
    assign _131 = _3295;
    always @(posedge _209) begin
        if (_223)
            _1039 <= _2929;
        else
            _1039 <= _131;
    end
    assign _1613 = { _3573,
                     _1039 };
    assign _1610 = { _3573,
                     _1035 };
    assign _1607 = { _3573,
                     _1317 };
    assign _1604 = { _3573,
                     _1603 };
    assign _1600 = { _3573,
                     _1599 };
    assign _1605 = _1600 + _1604;
    assign _1608 = _1605 + _1607;
    assign _1611 = _1608 + _1610;
    assign _1614 = _1611 + _1613;
    assign _1616 = _1614 < _3576;
    assign _1617 = _1321 & _1616;
    assign _3296 = ~ _1617;
    assign _3297 = _1321 & _3296;
    assign _3298 = _221 ? _3297 : _1321;
    assign _3299 = _531 ? _1317 : _3298;
    assign _132 = _3299;
    always @(posedge _209) begin
        if (_223)
            _1321 <= _2929;
        else
            _1321 <= _132;
    end
    assign _1346 = { _3573,
                     _1321 };
    assign _1343 = { _3573,
                     _1317 };
    assign _1341 = { _3573,
                     _1340 };
    assign _1344 = _1341 + _1343;
    assign _1347 = _1344 + _1346;
    assign _1350 = _1347 + _1349;
    assign _1353 = _1350 + _1352;
    assign _1356 = _1353 + _1355;
    assign _1359 = _1356 + _1358;
    assign _1362 = _1359 + _1361;
    assign _1364 = _1362 < _3576;
    assign _1365 = _1035 & _1364;
    assign _3300 = ~ _1365;
    assign _3301 = _1035 & _3300;
    assign _3302 = _221 ? _3301 : _1035;
    assign _3303 = _531 ? _1058 : _3302;
    assign _133 = _3303;
    always @(posedge _209) begin
        if (_223)
            _1035 <= _2929;
        else
            _1035 <= _133;
    end
    assign _1382 = { _3573,
                     _1035 };
    assign _1379 = { _3573,
                     _1088 };
    assign _1376 = { _3573,
                     _1317 };
    assign _1373 = { _3573,
                     _1340 };
    assign _1371 = { _3573,
                     _1370 };
    assign _1374 = _1371 + _1373;
    assign _1377 = _1374 + _1376;
    assign _1380 = _1377 + _1379;
    assign _1383 = _1380 + _1382;
    assign _1386 = _1383 + _1385;
    assign _1389 = _1386 + _1388;
    assign _1392 = _1389 + _1391;
    assign _1394 = _1392 < _3576;
    assign _1395 = _1058 & _1394;
    assign _3304 = ~ _1395;
    assign _3305 = _1058 & _3304;
    assign _3306 = _221 ? _3305 : _1058;
    assign _3307 = _531 ? _1088 : _3306;
    assign _134 = _3307;
    always @(posedge _209) begin
        if (_223)
            _1058 <= _2929;
        else
            _1058 <= _134;
    end
    assign _1412 = { _3573,
                     _1058 };
    assign _1409 = { _3573,
                     _1118 };
    assign _1406 = { _3573,
                     _1340 };
    assign _1403 = { _3573,
                     _1370 };
    assign _1401 = { _3573,
                     _1400 };
    assign _1404 = _1401 + _1403;
    assign _1407 = _1404 + _1406;
    assign _1410 = _1407 + _1409;
    assign _1413 = _1410 + _1412;
    assign _1416 = _1413 + _1415;
    assign _1419 = _1416 + _1418;
    assign _1422 = _1419 + _1421;
    assign _1424 = _1422 < _3576;
    assign _1425 = _1088 & _1424;
    assign _3308 = ~ _1425;
    assign _3309 = _1088 & _3308;
    assign _3310 = _221 ? _3309 : _1088;
    assign _3311 = _531 ? _1118 : _3310;
    assign _135 = _3311;
    always @(posedge _209) begin
        if (_223)
            _1088 <= _2929;
        else
            _1088 <= _135;
    end
    assign _1442 = { _3573,
                     _1088 };
    assign _1439 = { _3573,
                     _1148 };
    assign _1436 = { _3573,
                     _1370 };
    assign _1433 = { _3573,
                     _1400 };
    assign _1431 = { _3573,
                     _1430 };
    assign _1434 = _1431 + _1433;
    assign _1437 = _1434 + _1436;
    assign _1440 = _1437 + _1439;
    assign _1443 = _1440 + _1442;
    assign _1446 = _1443 + _1445;
    assign _1449 = _1446 + _1448;
    assign _1452 = _1449 + _1451;
    assign _1454 = _1452 < _3576;
    assign _1455 = _1118 & _1454;
    assign _3312 = ~ _1455;
    assign _3313 = _1118 & _3312;
    assign _3314 = _221 ? _3313 : _1118;
    assign _3315 = _531 ? _1148 : _3314;
    assign _136 = _3315;
    always @(posedge _209) begin
        if (_223)
            _1118 <= _2929;
        else
            _1118 <= _136;
    end
    assign _1472 = { _3573,
                     _1118 };
    assign _1469 = { _3573,
                     _1178 };
    assign _1466 = { _3573,
                     _1400 };
    assign _1463 = { _3573,
                     _1430 };
    assign _1461 = { _3573,
                     _1460 };
    assign _1464 = _1461 + _1463;
    assign _1467 = _1464 + _1466;
    assign _1470 = _1467 + _1469;
    assign _1473 = _1470 + _1472;
    assign _1476 = _1473 + _1475;
    assign _1479 = _1476 + _1478;
    assign _1482 = _1479 + _1481;
    assign _1484 = _1482 < _3576;
    assign _1485 = _1148 & _1484;
    assign _3316 = ~ _1485;
    assign _3317 = _1148 & _3316;
    assign _3318 = _221 ? _3317 : _1148;
    assign _3319 = _531 ? _1178 : _3318;
    assign _137 = _3319;
    always @(posedge _209) begin
        if (_223)
            _1148 <= _2929;
        else
            _1148 <= _137;
    end
    assign _1502 = { _3573,
                     _1148 };
    assign _1499 = { _3573,
                     _1208 };
    assign _1496 = { _3573,
                     _1430 };
    assign _1493 = { _3573,
                     _1460 };
    assign _1491 = { _3573,
                     _1490 };
    assign _1494 = _1491 + _1493;
    assign _1497 = _1494 + _1496;
    assign _1500 = _1497 + _1499;
    assign _1503 = _1500 + _1502;
    assign _1506 = _1503 + _1505;
    assign _1509 = _1506 + _1508;
    assign _1512 = _1509 + _1511;
    assign _1514 = _1512 < _3576;
    assign _1515 = _1178 & _1514;
    assign _3320 = ~ _1515;
    assign _3321 = _1178 & _3320;
    assign _3322 = _221 ? _3321 : _1178;
    assign _3323 = _531 ? _1208 : _3322;
    assign _138 = _3323;
    always @(posedge _209) begin
        if (_223)
            _1178 <= _2929;
        else
            _1178 <= _138;
    end
    assign _1532 = { _3573,
                     _1178 };
    assign _1529 = { _3573,
                     _1238 };
    assign _1526 = { _3573,
                     _1460 };
    assign _1523 = { _3573,
                     _1490 };
    assign _1521 = { _3573,
                     _1520 };
    assign _1524 = _1521 + _1523;
    assign _1527 = _1524 + _1526;
    assign _1530 = _1527 + _1529;
    assign _1533 = _1530 + _1532;
    assign _1536 = _1533 + _1535;
    assign _1539 = _1536 + _1538;
    assign _1542 = _1539 + _1541;
    assign _1544 = _1542 < _3576;
    assign _1545 = _1208 & _1544;
    assign _3324 = ~ _1545;
    assign _3325 = _1208 & _3324;
    assign _3326 = _221 ? _3325 : _1208;
    assign _3327 = _531 ? _1238 : _3326;
    assign _139 = _3327;
    always @(posedge _209) begin
        if (_223)
            _1208 <= _2929;
        else
            _1208 <= _139;
    end
    assign _1562 = { _3573,
                     _1208 };
    assign _1559 = { _3573,
                     _1268 };
    assign _1556 = { _3573,
                     _1490 };
    assign _1553 = { _3573,
                     _1520 };
    assign _1551 = { _3573,
                     _1550 };
    assign _1554 = _1551 + _1553;
    assign _1557 = _1554 + _1556;
    assign _1560 = _1557 + _1559;
    assign _1563 = _1560 + _1562;
    assign _1566 = _1563 + _1565;
    assign _1569 = _1566 + _1568;
    assign _1572 = _1569 + _1571;
    assign _1574 = _1572 < _3576;
    assign _1575 = _1238 & _1574;
    assign _3328 = ~ _1575;
    assign _3329 = _1238 & _3328;
    assign _3330 = _221 ? _3329 : _1238;
    assign _3331 = _531 ? _1268 : _3330;
    assign _140 = _3331;
    always @(posedge _209) begin
        if (_223)
            _1238 <= _2929;
        else
            _1238 <= _140;
    end
    assign _1584 = { _3573,
                     _1238 };
    assign _1581 = { _3573,
                     _1520 };
    assign _1579 = { _3573,
                     _1550 };
    assign _1582 = _1579 + _1581;
    assign _1585 = _1582 + _1584;
    assign _1588 = _1585 + _1587;
    assign _1591 = _1588 + _1590;
    assign _1593 = _1591 < _3576;
    assign _1594 = _1268 & _1593;
    assign _3332 = ~ _1594;
    assign _3333 = _1268 & _3332;
    assign _3334 = _221 ? _3333 : _1268;
    assign _3335 = _531 ? _1321 : _3334;
    assign _141 = _3335;
    always @(posedge _209) begin
        if (_223)
            _1268 <= _2929;
        else
            _1268 <= _141;
    end
    assign _1869 = { _3573,
                     _1268 };
    assign _1866 = { _3573,
                     _1520 };
    assign _1863 = { _3573,
                     _1802 };
    assign _1861 = { _3573,
                     _1832 };
    assign _1864 = _1861 + _1863;
    assign _1867 = _1864 + _1866;
    assign _1870 = _1867 + _1869;
    assign _1873 = _1870 + _1872;
    assign _1875 = _1873 < _3576;
    assign _1876 = _1550 & _1875;
    assign _3336 = ~ _1876;
    assign _3337 = _1550 & _3336;
    assign _3338 = _221 ? _3337 : _1550;
    assign _3339 = _531 ? _1603 : _3338;
    assign _142 = _3339;
    always @(posedge _209) begin
        if (_223)
            _1550 <= _2929;
        else
            _1550 <= _142;
    end
    assign _1841 = { _3573,
                     _1550 };
    assign _1838 = { _3573,
                     _1772 };
    assign _1835 = { _3573,
                     _1802 };
    assign _1833 = { _3573,
                     _1832 };
    assign _1836 = _1833 + _1835;
    assign _1839 = _1836 + _1838;
    assign _1842 = _1839 + _1841;
    assign _1845 = _1842 + _1844;
    assign _1848 = _1845 + _1847;
    assign _1851 = _1848 + _1850;
    assign _1854 = _1851 + _1853;
    assign _1856 = _1854 < _3576;
    assign _1857 = _1520 & _1856;
    assign _3340 = ~ _1857;
    assign _3341 = _1520 & _3340;
    assign _3342 = _221 ? _3341 : _1520;
    assign _3343 = _531 ? _1550 : _3342;
    assign _143 = _3343;
    always @(posedge _209) begin
        if (_223)
            _1520 <= _2929;
        else
            _1520 <= _143;
    end
    assign _1811 = { _3573,
                     _1520 };
    assign _1808 = { _3573,
                     _1742 };
    assign _1805 = { _3573,
                     _1772 };
    assign _1803 = { _3573,
                     _1802 };
    assign _1806 = _1803 + _1805;
    assign _1809 = _1806 + _1808;
    assign _1812 = _1809 + _1811;
    assign _1815 = _1812 + _1814;
    assign _1818 = _1815 + _1817;
    assign _1821 = _1818 + _1820;
    assign _1824 = _1821 + _1823;
    assign _1826 = _1824 < _3576;
    assign _1827 = _1490 & _1826;
    assign _3344 = ~ _1827;
    assign _3345 = _1490 & _3344;
    assign _3346 = _221 ? _3345 : _1490;
    assign _3347 = _531 ? _1520 : _3346;
    assign _144 = _3347;
    always @(posedge _209) begin
        if (_223)
            _1490 <= _2929;
        else
            _1490 <= _144;
    end
    assign _1781 = { _3573,
                     _1490 };
    assign _1778 = { _3573,
                     _1712 };
    assign _1775 = { _3573,
                     _1742 };
    assign _1773 = { _3573,
                     _1772 };
    assign _1776 = _1773 + _1775;
    assign _1779 = _1776 + _1778;
    assign _1782 = _1779 + _1781;
    assign _1785 = _1782 + _1784;
    assign _1788 = _1785 + _1787;
    assign _1791 = _1788 + _1790;
    assign _1794 = _1791 + _1793;
    assign _1796 = _1794 < _3576;
    assign _1797 = _1460 & _1796;
    assign _3348 = ~ _1797;
    assign _3349 = _1460 & _3348;
    assign _3350 = _221 ? _3349 : _1460;
    assign _3351 = _531 ? _1490 : _3350;
    assign _145 = _3351;
    always @(posedge _209) begin
        if (_223)
            _1460 <= _2929;
        else
            _1460 <= _145;
    end
    assign _1751 = { _3573,
                     _1460 };
    assign _1748 = { _3573,
                     _1682 };
    assign _1745 = { _3573,
                     _1712 };
    assign _1743 = { _3573,
                     _1742 };
    assign _1746 = _1743 + _1745;
    assign _1749 = _1746 + _1748;
    assign _1752 = _1749 + _1751;
    assign _1755 = _1752 + _1754;
    assign _1758 = _1755 + _1757;
    assign _1761 = _1758 + _1760;
    assign _1764 = _1761 + _1763;
    assign _1766 = _1764 < _3576;
    assign _1767 = _1430 & _1766;
    assign _3352 = ~ _1767;
    assign _3353 = _1430 & _3352;
    assign _3354 = _221 ? _3353 : _1430;
    assign _3355 = _531 ? _1460 : _3354;
    assign _146 = _3355;
    always @(posedge _209) begin
        if (_223)
            _1430 <= _2929;
        else
            _1430 <= _146;
    end
    assign _1721 = { _3573,
                     _1430 };
    assign _1718 = { _3573,
                     _1652 };
    assign _1715 = { _3573,
                     _1682 };
    assign _1713 = { _3573,
                     _1712 };
    assign _1716 = _1713 + _1715;
    assign _1719 = _1716 + _1718;
    assign _1722 = _1719 + _1721;
    assign _1725 = _1722 + _1724;
    assign _1728 = _1725 + _1727;
    assign _1731 = _1728 + _1730;
    assign _1734 = _1731 + _1733;
    assign _1736 = _1734 < _3576;
    assign _1737 = _1400 & _1736;
    assign _3356 = ~ _1737;
    assign _3357 = _1400 & _3356;
    assign _3358 = _221 ? _3357 : _1400;
    assign _3359 = _531 ? _1430 : _3358;
    assign _147 = _3359;
    always @(posedge _209) begin
        if (_223)
            _1400 <= _2929;
        else
            _1400 <= _147;
    end
    assign _1691 = { _3573,
                     _1400 };
    assign _1688 = { _3573,
                     _1622 };
    assign _1685 = { _3573,
                     _1652 };
    assign _1683 = { _3573,
                     _1682 };
    assign _1686 = _1683 + _1685;
    assign _1689 = _1686 + _1688;
    assign _1692 = _1689 + _1691;
    assign _1695 = _1692 + _1694;
    assign _1698 = _1695 + _1697;
    assign _1701 = _1698 + _1700;
    assign _1704 = _1701 + _1703;
    assign _1706 = _1704 < _3576;
    assign _1707 = _1370 & _1706;
    assign _3360 = ~ _1707;
    assign _3361 = _1370 & _3360;
    assign _3362 = _221 ? _3361 : _1370;
    assign _3363 = _531 ? _1400 : _3362;
    assign _148 = _3363;
    always @(posedge _209) begin
        if (_223)
            _1370 <= _2929;
        else
            _1370 <= _148;
    end
    assign _1661 = { _3573,
                     _1370 };
    assign _1658 = { _3573,
                     _1599 };
    assign _1655 = { _3573,
                     _1622 };
    assign _1653 = { _3573,
                     _1652 };
    assign _1656 = _1653 + _1655;
    assign _1659 = _1656 + _1658;
    assign _1662 = _1659 + _1661;
    assign _1665 = _1662 + _1664;
    assign _1668 = _1665 + _1667;
    assign _1671 = _1668 + _1670;
    assign _1674 = _1671 + _1673;
    assign _1676 = _1674 < _3576;
    assign _1677 = _1340 & _1676;
    assign _3364 = ~ _1677;
    assign _3365 = _1340 & _3364;
    assign _3366 = _221 ? _3365 : _1340;
    assign _3367 = _531 ? _1370 : _3366;
    assign _149 = _3367;
    always @(posedge _209) begin
        if (_223)
            _1340 <= _2929;
        else
            _1340 <= _149;
    end
    assign _1631 = { _3573,
                     _1340 };
    assign _1628 = { _3573,
                     _1603 };
    assign _1625 = { _3573,
                     _1599 };
    assign _1623 = { _3573,
                     _1622 };
    assign _1626 = _1623 + _1625;
    assign _1629 = _1626 + _1628;
    assign _1632 = _1629 + _1631;
    assign _1635 = _1632 + _1634;
    assign _1638 = _1635 + _1637;
    assign _1641 = _1638 + _1640;
    assign _1644 = _1641 + _1643;
    assign _1646 = _1644 < _3576;
    assign _1647 = _1317 & _1646;
    assign _3368 = ~ _1647;
    assign _3369 = _1317 & _3368;
    assign _3370 = _221 ? _3369 : _1317;
    assign _3371 = _531 ? _1340 : _3370;
    assign _150 = _3371;
    always @(posedge _209) begin
        if (_223)
            _1317 <= _2929;
        else
            _1317 <= _150;
    end
    assign _1892 = { _3573,
                     _1317 };
    assign _1889 = { _3573,
                     _1599 };
    assign _1886 = { _3573,
                     _1885 };
    assign _1882 = { _3573,
                     _1881 };
    assign _1887 = _1882 + _1886;
    assign _1890 = _1887 + _1889;
    assign _1893 = _1890 + _1892;
    assign _1896 = _1893 + _1895;
    assign _1898 = _1896 < _3576;
    assign _1899 = _1603 & _1898;
    assign _3372 = ~ _1899;
    assign _3373 = _1603 & _3372;
    assign _3374 = _221 ? _3373 : _1603;
    assign _3375 = _531 ? _1599 : _3374;
    assign _151 = _3375;
    always @(posedge _209) begin
        if (_223)
            _1603 <= _2929;
        else
            _1603 <= _151;
    end
    assign _2177 = { _3573,
                     _1603 };
    assign _2174 = { _3573,
                     _1599 };
    assign _2171 = { _3573,
                     _1881 };
    assign _2168 = { _3573,
                     _2167 };
    assign _2164 = { _3573,
                     _2163 };
    assign _2169 = _2164 + _2168;
    assign _2172 = _2169 + _2171;
    assign _2175 = _2172 + _2174;
    assign _2178 = _2175 + _2177;
    assign _2180 = _2178 < _3576;
    assign _2181 = _1885 & _2180;
    assign _3376 = ~ _2181;
    assign _3377 = _1885 & _3376;
    assign _3378 = _221 ? _3377 : _1885;
    assign _3379 = _531 ? _1881 : _3378;
    assign _152 = _3379;
    always @(posedge _209) begin
        if (_223)
            _1885 <= _2929;
        else
            _1885 <= _152;
    end
    assign _1910 = { _3573,
                     _1885 };
    assign _1907 = { _3573,
                     _1881 };
    assign _1905 = { _3573,
                     _1904 };
    assign _1908 = _1905 + _1907;
    assign _1911 = _1908 + _1910;
    assign _1914 = _1911 + _1913;
    assign _1917 = _1914 + _1916;
    assign _1920 = _1917 + _1919;
    assign _1923 = _1920 + _1922;
    assign _1926 = _1923 + _1925;
    assign _1928 = _1926 < _3576;
    assign _1929 = _1599 & _1928;
    assign _3380 = ~ _1929;
    assign _3381 = _1599 & _3380;
    assign _3382 = _221 ? _3381 : _1599;
    assign _3383 = _531 ? _1622 : _3382;
    assign _153 = _3383;
    always @(posedge _209) begin
        if (_223)
            _1599 <= _2929;
        else
            _1599 <= _153;
    end
    assign _1946 = { _3573,
                     _1599 };
    assign _1943 = { _3573,
                     _1652 };
    assign _1940 = { _3573,
                     _1881 };
    assign _1937 = { _3573,
                     _1904 };
    assign _1935 = { _3573,
                     _1934 };
    assign _1938 = _1935 + _1937;
    assign _1941 = _1938 + _1940;
    assign _1944 = _1941 + _1943;
    assign _1947 = _1944 + _1946;
    assign _1950 = _1947 + _1949;
    assign _1953 = _1950 + _1952;
    assign _1956 = _1953 + _1955;
    assign _1958 = _1956 < _3576;
    assign _1959 = _1622 & _1958;
    assign _3384 = ~ _1959;
    assign _3385 = _1622 & _3384;
    assign _3386 = _221 ? _3385 : _1622;
    assign _3387 = _531 ? _1652 : _3386;
    assign _154 = _3387;
    always @(posedge _209) begin
        if (_223)
            _1622 <= _2929;
        else
            _1622 <= _154;
    end
    assign _1976 = { _3573,
                     _1622 };
    assign _1973 = { _3573,
                     _1682 };
    assign _1970 = { _3573,
                     _1904 };
    assign _1967 = { _3573,
                     _1934 };
    assign _1965 = { _3573,
                     _1964 };
    assign _1968 = _1965 + _1967;
    assign _1971 = _1968 + _1970;
    assign _1974 = _1971 + _1973;
    assign _1977 = _1974 + _1976;
    assign _1980 = _1977 + _1979;
    assign _1983 = _1980 + _1982;
    assign _1986 = _1983 + _1985;
    assign _1988 = _1986 < _3576;
    assign _1989 = _1652 & _1988;
    assign _3388 = ~ _1989;
    assign _3389 = _1652 & _3388;
    assign _3390 = _221 ? _3389 : _1652;
    assign _3391 = _531 ? _1682 : _3390;
    assign _155 = _3391;
    always @(posedge _209) begin
        if (_223)
            _1652 <= _2929;
        else
            _1652 <= _155;
    end
    assign _2006 = { _3573,
                     _1652 };
    assign _2003 = { _3573,
                     _1712 };
    assign _2000 = { _3573,
                     _1934 };
    assign _1997 = { _3573,
                     _1964 };
    assign _1995 = { _3573,
                     _1994 };
    assign _1998 = _1995 + _1997;
    assign _2001 = _1998 + _2000;
    assign _2004 = _2001 + _2003;
    assign _2007 = _2004 + _2006;
    assign _2010 = _2007 + _2009;
    assign _2013 = _2010 + _2012;
    assign _2016 = _2013 + _2015;
    assign _2018 = _2016 < _3576;
    assign _2019 = _1682 & _2018;
    assign _3392 = ~ _2019;
    assign _3393 = _1682 & _3392;
    assign _3394 = _221 ? _3393 : _1682;
    assign _3395 = _531 ? _1712 : _3394;
    assign _156 = _3395;
    always @(posedge _209) begin
        if (_223)
            _1682 <= _2929;
        else
            _1682 <= _156;
    end
    assign _2036 = { _3573,
                     _1682 };
    assign _2033 = { _3573,
                     _1742 };
    assign _2030 = { _3573,
                     _1964 };
    assign _2027 = { _3573,
                     _1994 };
    assign _2025 = { _3573,
                     _2024 };
    assign _2028 = _2025 + _2027;
    assign _2031 = _2028 + _2030;
    assign _2034 = _2031 + _2033;
    assign _2037 = _2034 + _2036;
    assign _2040 = _2037 + _2039;
    assign _2043 = _2040 + _2042;
    assign _2046 = _2043 + _2045;
    assign _2048 = _2046 < _3576;
    assign _2049 = _1712 & _2048;
    assign _3396 = ~ _2049;
    assign _3397 = _1712 & _3396;
    assign _3398 = _221 ? _3397 : _1712;
    assign _3399 = _531 ? _1742 : _3398;
    assign _157 = _3399;
    always @(posedge _209) begin
        if (_223)
            _1712 <= _2929;
        else
            _1712 <= _157;
    end
    assign _2066 = { _3573,
                     _1712 };
    assign _2063 = { _3573,
                     _1772 };
    assign _2060 = { _3573,
                     _1994 };
    assign _2057 = { _3573,
                     _2024 };
    assign _2055 = { _3573,
                     _2054 };
    assign _2058 = _2055 + _2057;
    assign _2061 = _2058 + _2060;
    assign _2064 = _2061 + _2063;
    assign _2067 = _2064 + _2066;
    assign _2070 = _2067 + _2069;
    assign _2073 = _2070 + _2072;
    assign _2076 = _2073 + _2075;
    assign _2078 = _2076 < _3576;
    assign _2079 = _1742 & _2078;
    assign _3400 = ~ _2079;
    assign _3401 = _1742 & _3400;
    assign _3402 = _221 ? _3401 : _1742;
    assign _3403 = _531 ? _1772 : _3402;
    assign _158 = _3403;
    always @(posedge _209) begin
        if (_223)
            _1742 <= _2929;
        else
            _1742 <= _158;
    end
    assign _2096 = { _3573,
                     _1742 };
    assign _2093 = { _3573,
                     _1802 };
    assign _2090 = { _3573,
                     _2024 };
    assign _2087 = { _3573,
                     _2054 };
    assign _2085 = { _3573,
                     _2084 };
    assign _2088 = _2085 + _2087;
    assign _2091 = _2088 + _2090;
    assign _2094 = _2091 + _2093;
    assign _2097 = _2094 + _2096;
    assign _2100 = _2097 + _2099;
    assign _2103 = _2100 + _2102;
    assign _2106 = _2103 + _2105;
    assign _2108 = _2106 < _3576;
    assign _2109 = _1772 & _2108;
    assign _3404 = ~ _2109;
    assign _3405 = _1772 & _3404;
    assign _3406 = _221 ? _3405 : _1772;
    assign _3407 = _531 ? _1802 : _3406;
    assign _159 = _3407;
    always @(posedge _209) begin
        if (_223)
            _1772 <= _2929;
        else
            _1772 <= _159;
    end
    assign _2126 = { _3573,
                     _1772 };
    assign _2123 = { _3573,
                     _1832 };
    assign _2120 = { _3573,
                     _2054 };
    assign _2117 = { _3573,
                     _2084 };
    assign _2115 = { _3573,
                     _2114 };
    assign _2118 = _2115 + _2117;
    assign _2121 = _2118 + _2120;
    assign _2124 = _2121 + _2123;
    assign _2127 = _2124 + _2126;
    assign _2130 = _2127 + _2129;
    assign _2133 = _2130 + _2132;
    assign _2136 = _2133 + _2135;
    assign _2138 = _2136 < _3576;
    assign _2139 = _1802 & _2138;
    assign _3408 = ~ _2139;
    assign _3409 = _1802 & _3408;
    assign _3410 = _221 ? _3409 : _1802;
    assign _3411 = _531 ? _1832 : _3410;
    assign _160 = _3411;
    always @(posedge _209) begin
        if (_223)
            _1802 <= _2929;
        else
            _1802 <= _160;
    end
    assign _2148 = { _3573,
                     _1802 };
    assign _2145 = { _3573,
                     _2084 };
    assign _2143 = { _3573,
                     _2114 };
    assign _2146 = _2143 + _2145;
    assign _2149 = _2146 + _2148;
    assign _2152 = _2149 + _2151;
    assign _2155 = _2152 + _2154;
    assign _2157 = _2155 < _3576;
    assign _2158 = _1832 & _2157;
    assign _3412 = ~ _2158;
    assign _3413 = _1832 & _3412;
    assign _3414 = _221 ? _3413 : _1832;
    assign _3415 = _531 ? _1885 : _3414;
    assign _161 = _3415;
    always @(posedge _209) begin
        if (_223)
            _1832 <= _2929;
        else
            _1832 <= _161;
    end
    assign _2433 = { _3573,
                     _1832 };
    assign _2430 = { _3573,
                     _2084 };
    assign _2427 = { _3573,
                     _2366 };
    assign _2425 = { _3573,
                     _2396 };
    assign _2428 = _2425 + _2427;
    assign _2431 = _2428 + _2430;
    assign _2434 = _2431 + _2433;
    assign _2437 = _2434 + _2436;
    assign _2439 = _2437 < _3576;
    assign _2440 = _2114 & _2439;
    assign _3416 = ~ _2440;
    assign _3417 = _2114 & _3416;
    assign _3418 = _221 ? _3417 : _2114;
    assign _3419 = _531 ? _2167 : _3418;
    assign _162 = _3419;
    always @(posedge _209) begin
        if (_223)
            _2114 <= _2929;
        else
            _2114 <= _162;
    end
    assign _2405 = { _3573,
                     _2114 };
    assign _2402 = { _3573,
                     _2336 };
    assign _2399 = { _3573,
                     _2366 };
    assign _2397 = { _3573,
                     _2396 };
    assign _2400 = _2397 + _2399;
    assign _2403 = _2400 + _2402;
    assign _2406 = _2403 + _2405;
    assign _2409 = _2406 + _2408;
    assign _2412 = _2409 + _2411;
    assign _2415 = _2412 + _2414;
    assign _2418 = _2415 + _2417;
    assign _2420 = _2418 < _3576;
    assign _2421 = _2084 & _2420;
    assign _3420 = ~ _2421;
    assign _3421 = _2084 & _3420;
    assign _3422 = _221 ? _3421 : _2084;
    assign _3423 = _531 ? _2114 : _3422;
    assign _163 = _3423;
    always @(posedge _209) begin
        if (_223)
            _2084 <= _2929;
        else
            _2084 <= _163;
    end
    assign _2375 = { _3573,
                     _2084 };
    assign _2372 = { _3573,
                     _2306 };
    assign _2369 = { _3573,
                     _2336 };
    assign _2367 = { _3573,
                     _2366 };
    assign _2370 = _2367 + _2369;
    assign _2373 = _2370 + _2372;
    assign _2376 = _2373 + _2375;
    assign _2379 = _2376 + _2378;
    assign _2382 = _2379 + _2381;
    assign _2385 = _2382 + _2384;
    assign _2388 = _2385 + _2387;
    assign _2390 = _2388 < _3576;
    assign _2391 = _2054 & _2390;
    assign _3424 = ~ _2391;
    assign _3425 = _2054 & _3424;
    assign _3426 = _221 ? _3425 : _2054;
    assign _3427 = _531 ? _2084 : _3426;
    assign _164 = _3427;
    always @(posedge _209) begin
        if (_223)
            _2054 <= _2929;
        else
            _2054 <= _164;
    end
    assign _2345 = { _3573,
                     _2054 };
    assign _2342 = { _3573,
                     _2276 };
    assign _2339 = { _3573,
                     _2306 };
    assign _2337 = { _3573,
                     _2336 };
    assign _2340 = _2337 + _2339;
    assign _2343 = _2340 + _2342;
    assign _2346 = _2343 + _2345;
    assign _2349 = _2346 + _2348;
    assign _2352 = _2349 + _2351;
    assign _2355 = _2352 + _2354;
    assign _2358 = _2355 + _2357;
    assign _2360 = _2358 < _3576;
    assign _2361 = _2024 & _2360;
    assign _3428 = ~ _2361;
    assign _3429 = _2024 & _3428;
    assign _3430 = _221 ? _3429 : _2024;
    assign _3431 = _531 ? _2054 : _3430;
    assign _165 = _3431;
    always @(posedge _209) begin
        if (_223)
            _2024 <= _2929;
        else
            _2024 <= _165;
    end
    assign _2315 = { _3573,
                     _2024 };
    assign _2312 = { _3573,
                     _2246 };
    assign _2309 = { _3573,
                     _2276 };
    assign _2307 = { _3573,
                     _2306 };
    assign _2310 = _2307 + _2309;
    assign _2313 = _2310 + _2312;
    assign _2316 = _2313 + _2315;
    assign _2319 = _2316 + _2318;
    assign _2322 = _2319 + _2321;
    assign _2325 = _2322 + _2324;
    assign _2328 = _2325 + _2327;
    assign _2330 = _2328 < _3576;
    assign _2331 = _1994 & _2330;
    assign _3432 = ~ _2331;
    assign _3433 = _1994 & _3432;
    assign _3434 = _221 ? _3433 : _1994;
    assign _3435 = _531 ? _2024 : _3434;
    assign _166 = _3435;
    always @(posedge _209) begin
        if (_223)
            _1994 <= _2929;
        else
            _1994 <= _166;
    end
    assign _2285 = { _3573,
                     _1994 };
    assign _2282 = { _3573,
                     _2216 };
    assign _2279 = { _3573,
                     _2246 };
    assign _2277 = { _3573,
                     _2276 };
    assign _2280 = _2277 + _2279;
    assign _2283 = _2280 + _2282;
    assign _2286 = _2283 + _2285;
    assign _2289 = _2286 + _2288;
    assign _2292 = _2289 + _2291;
    assign _2295 = _2292 + _2294;
    assign _2298 = _2295 + _2297;
    assign _2300 = _2298 < _3576;
    assign _2301 = _1964 & _2300;
    assign _3436 = ~ _2301;
    assign _3437 = _1964 & _3436;
    assign _3438 = _221 ? _3437 : _1964;
    assign _3439 = _531 ? _1994 : _3438;
    assign _167 = _3439;
    always @(posedge _209) begin
        if (_223)
            _1964 <= _2929;
        else
            _1964 <= _167;
    end
    assign _2255 = { _3573,
                     _1964 };
    assign _2252 = { _3573,
                     _2186 };
    assign _2249 = { _3573,
                     _2216 };
    assign _2247 = { _3573,
                     _2246 };
    assign _2250 = _2247 + _2249;
    assign _2253 = _2250 + _2252;
    assign _2256 = _2253 + _2255;
    assign _2259 = _2256 + _2258;
    assign _2262 = _2259 + _2261;
    assign _2265 = _2262 + _2264;
    assign _2268 = _2265 + _2267;
    assign _2270 = _2268 < _3576;
    assign _2271 = _1934 & _2270;
    assign _3440 = ~ _2271;
    assign _3441 = _1934 & _3440;
    assign _3442 = _221 ? _3441 : _1934;
    assign _3443 = _531 ? _1964 : _3442;
    assign _168 = _3443;
    always @(posedge _209) begin
        if (_223)
            _1934 <= _2929;
        else
            _1934 <= _168;
    end
    assign _2225 = { _3573,
                     _1934 };
    assign _2222 = { _3573,
                     _2163 };
    assign _2219 = { _3573,
                     _2186 };
    assign _2217 = { _3573,
                     _2216 };
    assign _2220 = _2217 + _2219;
    assign _2223 = _2220 + _2222;
    assign _2226 = _2223 + _2225;
    assign _2229 = _2226 + _2228;
    assign _2232 = _2229 + _2231;
    assign _2235 = _2232 + _2234;
    assign _2238 = _2235 + _2237;
    assign _2240 = _2238 < _3576;
    assign _2241 = _1904 & _2240;
    assign _3444 = ~ _2241;
    assign _3445 = _1904 & _3444;
    assign _3446 = _221 ? _3445 : _1904;
    assign _3447 = _531 ? _1934 : _3446;
    assign _169 = _3447;
    always @(posedge _209) begin
        if (_223)
            _1904 <= _2929;
        else
            _1904 <= _169;
    end
    assign _2195 = { _3573,
                     _1904 };
    assign _2192 = { _3573,
                     _2167 };
    assign _2189 = { _3573,
                     _2163 };
    assign _2187 = { _3573,
                     _2186 };
    assign _2190 = _2187 + _2189;
    assign _2193 = _2190 + _2192;
    assign _2196 = _2193 + _2195;
    assign _2199 = _2196 + _2198;
    assign _2202 = _2199 + _2201;
    assign _2205 = _2202 + _2204;
    assign _2208 = _2205 + _2207;
    assign _2210 = _2208 < _3576;
    assign _2211 = _1881 & _2210;
    assign _3448 = ~ _2211;
    assign _3449 = _1881 & _3448;
    assign _3450 = _221 ? _3449 : _1881;
    assign _3451 = _531 ? _1904 : _3450;
    assign _170 = _3451;
    always @(posedge _209) begin
        if (_223)
            _1881 <= _2929;
        else
            _1881 <= _170;
    end
    assign _2456 = { _3573,
                     _1881 };
    assign _2453 = { _3573,
                     _2163 };
    assign _2450 = { _3573,
                     _2449 };
    assign _2446 = { _3573,
                     _2445 };
    assign _2451 = _2446 + _2450;
    assign _2454 = _2451 + _2453;
    assign _2457 = _2454 + _2456;
    assign _2460 = _2457 + _2459;
    assign _2462 = _2460 < _3576;
    assign _2463 = _2167 & _2462;
    assign _3452 = ~ _2463;
    assign _3453 = _2167 & _3452;
    assign _3454 = _221 ? _3453 : _2167;
    assign _3455 = _531 ? _2163 : _3454;
    assign _171 = _3455;
    always @(posedge _209) begin
        if (_223)
            _2167 <= _2929;
        else
            _2167 <= _171;
    end
    assign _2741 = { _3573,
                     _2167 };
    assign _2738 = { _3573,
                     _2163 };
    assign _2735 = { _3573,
                     _2445 };
    assign _2732 = { _3573,
                     _2731 };
    assign _2728 = { _3573,
                     _2727 };
    assign _2733 = _2728 + _2732;
    assign _2736 = _2733 + _2735;
    assign _2739 = _2736 + _2738;
    assign _2742 = _2739 + _2741;
    assign _2744 = _2742 < _3576;
    assign _2745 = _2449 & _2744;
    assign _3456 = ~ _2745;
    assign _3457 = _2449 & _3456;
    assign _3458 = _221 ? _3457 : _2449;
    assign _3459 = _531 ? _2445 : _3458;
    assign _172 = _3459;
    always @(posedge _209) begin
        if (_223)
            _2449 <= _2929;
        else
            _2449 <= _172;
    end
    assign _2474 = { _3573,
                     _2449 };
    assign _2471 = { _3573,
                     _2445 };
    assign _2469 = { _3573,
                     _2468 };
    assign _2472 = _2469 + _2471;
    assign _2475 = _2472 + _2474;
    assign _2478 = _2475 + _2477;
    assign _2481 = _2478 + _2480;
    assign _2484 = _2481 + _2483;
    assign _2487 = _2484 + _2486;
    assign _2490 = _2487 + _2489;
    assign _2492 = _2490 < _3576;
    assign _2493 = _2163 & _2492;
    assign _3460 = ~ _2493;
    assign _3461 = _2163 & _3460;
    assign _3462 = _221 ? _3461 : _2163;
    assign _3463 = _531 ? _2186 : _3462;
    assign _173 = _3463;
    always @(posedge _209) begin
        if (_223)
            _2163 <= _2929;
        else
            _2163 <= _173;
    end
    assign _2510 = { _3573,
                     _2163 };
    assign _2507 = { _3573,
                     _2216 };
    assign _2504 = { _3573,
                     _2445 };
    assign _2501 = { _3573,
                     _2468 };
    assign _2499 = { _3573,
                     _2498 };
    assign _2502 = _2499 + _2501;
    assign _2505 = _2502 + _2504;
    assign _2508 = _2505 + _2507;
    assign _2511 = _2508 + _2510;
    assign _2514 = _2511 + _2513;
    assign _2517 = _2514 + _2516;
    assign _2520 = _2517 + _2519;
    assign _2522 = _2520 < _3576;
    assign _2523 = _2186 & _2522;
    assign _3464 = ~ _2523;
    assign _3465 = _2186 & _3464;
    assign _3466 = _221 ? _3465 : _2186;
    assign _3467 = _531 ? _2216 : _3466;
    assign _174 = _3467;
    always @(posedge _209) begin
        if (_223)
            _2186 <= _2929;
        else
            _2186 <= _174;
    end
    assign _2540 = { _3573,
                     _2186 };
    assign _2537 = { _3573,
                     _2246 };
    assign _2534 = { _3573,
                     _2468 };
    assign _2531 = { _3573,
                     _2498 };
    assign _2529 = { _3573,
                     _2528 };
    assign _2532 = _2529 + _2531;
    assign _2535 = _2532 + _2534;
    assign _2538 = _2535 + _2537;
    assign _2541 = _2538 + _2540;
    assign _2544 = _2541 + _2543;
    assign _2547 = _2544 + _2546;
    assign _2550 = _2547 + _2549;
    assign _2552 = _2550 < _3576;
    assign _2553 = _2216 & _2552;
    assign _3468 = ~ _2553;
    assign _3469 = _2216 & _3468;
    assign _3470 = _221 ? _3469 : _2216;
    assign _3471 = _531 ? _2246 : _3470;
    assign _175 = _3471;
    always @(posedge _209) begin
        if (_223)
            _2216 <= _2929;
        else
            _2216 <= _175;
    end
    assign _2570 = { _3573,
                     _2216 };
    assign _2567 = { _3573,
                     _2276 };
    assign _2564 = { _3573,
                     _2498 };
    assign _2561 = { _3573,
                     _2528 };
    assign _2559 = { _3573,
                     _2558 };
    assign _2562 = _2559 + _2561;
    assign _2565 = _2562 + _2564;
    assign _2568 = _2565 + _2567;
    assign _2571 = _2568 + _2570;
    assign _2574 = _2571 + _2573;
    assign _2577 = _2574 + _2576;
    assign _2580 = _2577 + _2579;
    assign _2582 = _2580 < _3576;
    assign _2583 = _2246 & _2582;
    assign _3472 = ~ _2583;
    assign _3473 = _2246 & _3472;
    assign _3474 = _221 ? _3473 : _2246;
    assign _3475 = _531 ? _2276 : _3474;
    assign _176 = _3475;
    always @(posedge _209) begin
        if (_223)
            _2246 <= _2929;
        else
            _2246 <= _176;
    end
    assign _2600 = { _3573,
                     _2246 };
    assign _2597 = { _3573,
                     _2306 };
    assign _2594 = { _3573,
                     _2528 };
    assign _2591 = { _3573,
                     _2558 };
    assign _2589 = { _3573,
                     _2588 };
    assign _2592 = _2589 + _2591;
    assign _2595 = _2592 + _2594;
    assign _2598 = _2595 + _2597;
    assign _2601 = _2598 + _2600;
    assign _2604 = _2601 + _2603;
    assign _2607 = _2604 + _2606;
    assign _2610 = _2607 + _2609;
    assign _2612 = _2610 < _3576;
    assign _2613 = _2276 & _2612;
    assign _3476 = ~ _2613;
    assign _3477 = _2276 & _3476;
    assign _3478 = _221 ? _3477 : _2276;
    assign _3479 = _531 ? _2306 : _3478;
    assign _177 = _3479;
    always @(posedge _209) begin
        if (_223)
            _2276 <= _2929;
        else
            _2276 <= _177;
    end
    assign _2630 = { _3573,
                     _2276 };
    assign _2627 = { _3573,
                     _2336 };
    assign _2624 = { _3573,
                     _2558 };
    assign _2621 = { _3573,
                     _2588 };
    assign _2619 = { _3573,
                     _2618 };
    assign _2622 = _2619 + _2621;
    assign _2625 = _2622 + _2624;
    assign _2628 = _2625 + _2627;
    assign _2631 = _2628 + _2630;
    assign _2634 = _2631 + _2633;
    assign _2637 = _2634 + _2636;
    assign _2640 = _2637 + _2639;
    assign _2642 = _2640 < _3576;
    assign _2643 = _2306 & _2642;
    assign _3480 = ~ _2643;
    assign _3481 = _2306 & _3480;
    assign _3482 = _221 ? _3481 : _2306;
    assign _3483 = _531 ? _2336 : _3482;
    assign _178 = _3483;
    always @(posedge _209) begin
        if (_223)
            _2306 <= _2929;
        else
            _2306 <= _178;
    end
    assign _2660 = { _3573,
                     _2306 };
    assign _2657 = { _3573,
                     _2366 };
    assign _2654 = { _3573,
                     _2588 };
    assign _2651 = { _3573,
                     _2618 };
    assign _2649 = { _3573,
                     _2648 };
    assign _2652 = _2649 + _2651;
    assign _2655 = _2652 + _2654;
    assign _2658 = _2655 + _2657;
    assign _2661 = _2658 + _2660;
    assign _2664 = _2661 + _2663;
    assign _2667 = _2664 + _2666;
    assign _2670 = _2667 + _2669;
    assign _2672 = _2670 < _3576;
    assign _2673 = _2336 & _2672;
    assign _3484 = ~ _2673;
    assign _3485 = _2336 & _3484;
    assign _3486 = _221 ? _3485 : _2336;
    assign _3487 = _531 ? _2366 : _3486;
    assign _179 = _3487;
    always @(posedge _209) begin
        if (_223)
            _2336 <= _2929;
        else
            _2336 <= _179;
    end
    assign _2690 = { _3573,
                     _2336 };
    assign _2687 = { _3573,
                     _2396 };
    assign _2684 = { _3573,
                     _2618 };
    assign _2681 = { _3573,
                     _2648 };
    assign _2679 = { _3573,
                     _2678 };
    assign _2682 = _2679 + _2681;
    assign _2685 = _2682 + _2684;
    assign _2688 = _2685 + _2687;
    assign _2691 = _2688 + _2690;
    assign _2694 = _2691 + _2693;
    assign _2697 = _2694 + _2696;
    assign _2700 = _2697 + _2699;
    assign _2702 = _2700 < _3576;
    assign _2703 = _2366 & _2702;
    assign _3488 = ~ _2703;
    assign _3489 = _2366 & _3488;
    assign _3490 = _221 ? _3489 : _2366;
    assign _3491 = _531 ? _2396 : _3490;
    assign _180 = _3491;
    always @(posedge _209) begin
        if (_223)
            _2366 <= _2929;
        else
            _2366 <= _180;
    end
    assign _2712 = { _3573,
                     _2366 };
    assign _2709 = { _3573,
                     _2648 };
    assign _2707 = { _3573,
                     _2678 };
    assign _2710 = _2707 + _2709;
    assign _2713 = _2710 + _2712;
    assign _2716 = _2713 + _2715;
    assign _2719 = _2716 + _2718;
    assign _2721 = _2719 < _3576;
    assign _2722 = _2396 & _2721;
    assign _3492 = ~ _2722;
    assign _3493 = _2396 & _3492;
    assign _3494 = _221 ? _3493 : _2396;
    assign _3495 = _531 ? _2449 : _3494;
    assign _181 = _3495;
    always @(posedge _209) begin
        if (_223)
            _2396 <= _2929;
        else
            _2396 <= _181;
    end
    assign _2997 = { _3573,
                     _2396 };
    assign _2994 = { _3573,
                     _2648 };
    assign _2991 = { _3573,
                     _2930 };
    assign _2989 = { _3573,
                     _2960 };
    assign _2992 = _2989 + _2991;
    assign _2995 = _2992 + _2994;
    assign _2998 = _2995 + _2997;
    assign _3001 = _2998 + _3000;
    assign _3003 = _3001 < _3576;
    assign _3004 = _2678 & _3003;
    assign _3496 = ~ _3004;
    assign _3497 = _2678 & _3496;
    assign _3498 = _221 ? _3497 : _2678;
    assign _3499 = _531 ? _2731 : _3498;
    assign _182 = _3499;
    always @(posedge _209) begin
        if (_223)
            _2678 <= _2929;
        else
            _2678 <= _182;
    end
    assign _2969 = { _3573,
                     _2678 };
    assign _2966 = { _3573,
                     _2900 };
    assign _2963 = { _3573,
                     _2930 };
    assign _2961 = { _3573,
                     _2960 };
    assign _2964 = _2961 + _2963;
    assign _2967 = _2964 + _2966;
    assign _2970 = _2967 + _2969;
    assign _2973 = _2970 + _2972;
    assign _2976 = _2973 + _2975;
    assign _2979 = _2976 + _2978;
    assign _2982 = _2979 + _2981;
    assign _2984 = _2982 < _3576;
    assign _2985 = _2648 & _2984;
    assign _3500 = ~ _2985;
    assign _3501 = _2648 & _3500;
    assign _3502 = _221 ? _3501 : _2648;
    assign _3503 = _531 ? _2678 : _3502;
    assign _183 = _3503;
    always @(posedge _209) begin
        if (_223)
            _2648 <= _2929;
        else
            _2648 <= _183;
    end
    assign _2939 = { _3573,
                     _2648 };
    assign _2936 = { _3573,
                     _2870 };
    assign _2933 = { _3573,
                     _2900 };
    assign _2931 = { _3573,
                     _2930 };
    assign _2934 = _2931 + _2933;
    assign _2937 = _2934 + _2936;
    assign _2940 = _2937 + _2939;
    assign _2943 = _2940 + _2942;
    assign _2946 = _2943 + _2945;
    assign _2949 = _2946 + _2948;
    assign _2952 = _2949 + _2951;
    assign _2954 = _2952 < _3576;
    assign _2955 = _2618 & _2954;
    assign _3504 = ~ _2955;
    assign _3505 = _2618 & _3504;
    assign _3506 = _221 ? _3505 : _2618;
    assign _3507 = _531 ? _2648 : _3506;
    assign _184 = _3507;
    always @(posedge _209) begin
        if (_223)
            _2618 <= _2929;
        else
            _2618 <= _184;
    end
    assign _2909 = { _3573,
                     _2618 };
    assign _2906 = { _3573,
                     _2840 };
    assign _2903 = { _3573,
                     _2870 };
    assign _2901 = { _3573,
                     _2900 };
    assign _2904 = _2901 + _2903;
    assign _2907 = _2904 + _2906;
    assign _2910 = _2907 + _2909;
    assign _2913 = _2910 + _2912;
    assign _2916 = _2913 + _2915;
    assign _2919 = _2916 + _2918;
    assign _2922 = _2919 + _2921;
    assign _2924 = _2922 < _3576;
    assign _2925 = _2588 & _2924;
    assign _3508 = ~ _2925;
    assign _3509 = _2588 & _3508;
    assign _3510 = _221 ? _3509 : _2588;
    assign _3511 = _531 ? _2618 : _3510;
    assign _185 = _3511;
    always @(posedge _209) begin
        if (_223)
            _2588 <= _2929;
        else
            _2588 <= _185;
    end
    assign _2879 = { _3573,
                     _2588 };
    assign _2876 = { _3573,
                     _2810 };
    assign _2873 = { _3573,
                     _2840 };
    assign _2871 = { _3573,
                     _2870 };
    assign _2874 = _2871 + _2873;
    assign _2877 = _2874 + _2876;
    assign _2880 = _2877 + _2879;
    assign _2883 = _2880 + _2882;
    assign _2886 = _2883 + _2885;
    assign _2889 = _2886 + _2888;
    assign _2892 = _2889 + _2891;
    assign _2894 = _2892 < _3576;
    assign _2895 = _2558 & _2894;
    assign _3512 = ~ _2895;
    assign _3513 = _2558 & _3512;
    assign _3514 = _221 ? _3513 : _2558;
    assign _3515 = _531 ? _2588 : _3514;
    assign _186 = _3515;
    always @(posedge _209) begin
        if (_223)
            _2558 <= _2929;
        else
            _2558 <= _186;
    end
    assign _2849 = { _3573,
                     _2558 };
    assign _2846 = { _3573,
                     _2780 };
    assign _2843 = { _3573,
                     _2810 };
    assign _2841 = { _3573,
                     _2840 };
    assign _2844 = _2841 + _2843;
    assign _2847 = _2844 + _2846;
    assign _2850 = _2847 + _2849;
    assign _2853 = _2850 + _2852;
    assign _2856 = _2853 + _2855;
    assign _2859 = _2856 + _2858;
    assign _2862 = _2859 + _2861;
    assign _2864 = _2862 < _3576;
    assign _2865 = _2528 & _2864;
    assign _3516 = ~ _2865;
    assign _3517 = _2528 & _3516;
    assign _3518 = _221 ? _3517 : _2528;
    assign _3519 = _531 ? _2558 : _3518;
    assign _187 = _3519;
    always @(posedge _209) begin
        if (_223)
            _2528 <= _2929;
        else
            _2528 <= _187;
    end
    assign _2819 = { _3573,
                     _2528 };
    assign _2816 = { _3573,
                     _2750 };
    assign _2813 = { _3573,
                     _2780 };
    assign _2811 = { _3573,
                     _2810 };
    assign _2814 = _2811 + _2813;
    assign _2817 = _2814 + _2816;
    assign _2820 = _2817 + _2819;
    assign _2823 = _2820 + _2822;
    assign _2826 = _2823 + _2825;
    assign _2829 = _2826 + _2828;
    assign _2832 = _2829 + _2831;
    assign _2834 = _2832 < _3576;
    assign _2835 = _2498 & _2834;
    assign _3520 = ~ _2835;
    assign _3521 = _2498 & _3520;
    assign _3522 = _221 ? _3521 : _2498;
    assign _3523 = _531 ? _2528 : _3522;
    assign _188 = _3523;
    always @(posedge _209) begin
        if (_223)
            _2498 <= _2929;
        else
            _2498 <= _188;
    end
    assign _2789 = { _3573,
                     _2498 };
    assign _2786 = { _3573,
                     _2727 };
    assign _2783 = { _3573,
                     _2750 };
    assign _2781 = { _3573,
                     _2780 };
    assign _2784 = _2781 + _2783;
    assign _2787 = _2784 + _2786;
    assign _2790 = _2787 + _2789;
    assign _2793 = _2790 + _2792;
    assign _2796 = _2793 + _2795;
    assign _2799 = _2796 + _2798;
    assign _2802 = _2799 + _2801;
    assign _2804 = _2802 < _3576;
    assign _2805 = _2468 & _2804;
    assign _3524 = ~ _2805;
    assign _3525 = _2468 & _3524;
    assign _3526 = _221 ? _3525 : _2468;
    assign _3527 = _531 ? _2498 : _3526;
    assign _189 = _3527;
    always @(posedge _209) begin
        if (_223)
            _2468 <= _2929;
        else
            _2468 <= _189;
    end
    assign _2759 = { _3573,
                     _2468 };
    assign _2756 = { _3573,
                     _2731 };
    assign _2753 = { _3573,
                     _2727 };
    assign _2751 = { _3573,
                     _2750 };
    assign _2754 = _2751 + _2753;
    assign _2757 = _2754 + _2756;
    assign _2760 = _2757 + _2759;
    assign _2763 = _2760 + _2762;
    assign _2766 = _2763 + _2765;
    assign _2769 = _2766 + _2768;
    assign _2772 = _2769 + _2771;
    assign _2774 = _2772 < _3576;
    assign _2775 = _2445 & _2774;
    assign _3528 = ~ _2775;
    assign _3529 = _2445 & _3528;
    assign _3530 = _221 ? _3529 : _2445;
    assign _3531 = _531 ? _2468 : _3530;
    assign _190 = _3531;
    always @(posedge _209) begin
        if (_223)
            _2445 <= _2929;
        else
            _2445 <= _190;
    end
    assign _3010 = { _3573,
                     _2445 };
    assign _3008 = { _3573,
                     _2727 };
    assign _3011 = _3008 + _3010;
    assign _3014 = _3011 + _3013;
    assign _3016 = _3014 < _3576;
    assign _3017 = _2731 & _3016;
    assign _3532 = ~ _3017;
    assign _3533 = _2731 & _3532;
    assign _3534 = _221 ? _3533 : _2731;
    assign _3535 = _531 ? _2727 : _3534;
    assign _191 = _3535;
    always @(posedge _209) begin
        if (_223)
            _2731 <= _2929;
        else
            _2731 <= _191;
    end
    assign _3023 = { _3573,
                     _2731 };
    assign _3021 = { _3573,
                     _2750 };
    assign _3024 = _3021 + _3023;
    assign _3027 = _3024 + _3026;
    assign _3030 = _3027 + _3029;
    assign _3033 = _3030 + _3032;
    assign _3035 = _3033 < _3576;
    assign _3036 = _2727 & _3035;
    assign _3536 = ~ _3036;
    assign _3537 = _2727 & _3536;
    assign _3538 = _221 ? _3537 : _2727;
    assign _3539 = _531 ? _2750 : _3538;
    assign _192 = _3539;
    always @(posedge _209) begin
        if (_223)
            _2727 <= _2929;
        else
            _2727 <= _192;
    end
    assign _3042 = { _3573,
                     _2727 };
    assign _3040 = { _3573,
                     _2780 };
    assign _3043 = _3040 + _3042;
    assign _3046 = _3043 + _3045;
    assign _3049 = _3046 + _3048;
    assign _3052 = _3049 + _3051;
    assign _3054 = _3052 < _3576;
    assign _3055 = _2750 & _3054;
    assign _3540 = ~ _3055;
    assign _3541 = _2750 & _3540;
    assign _3542 = _221 ? _3541 : _2750;
    assign _3543 = _531 ? _2780 : _3542;
    assign _193 = _3543;
    always @(posedge _209) begin
        if (_223)
            _2750 <= _2929;
        else
            _2750 <= _193;
    end
    assign _3061 = { _3573,
                     _2750 };
    assign _3059 = { _3573,
                     _2810 };
    assign _3062 = _3059 + _3061;
    assign _3065 = _3062 + _3064;
    assign _3068 = _3065 + _3067;
    assign _3071 = _3068 + _3070;
    assign _3073 = _3071 < _3576;
    assign _3074 = _2780 & _3073;
    assign _3544 = ~ _3074;
    assign _3545 = _2780 & _3544;
    assign _3546 = _221 ? _3545 : _2780;
    assign _3547 = _531 ? _2810 : _3546;
    assign _194 = _3547;
    always @(posedge _209) begin
        if (_223)
            _2780 <= _2929;
        else
            _2780 <= _194;
    end
    assign _3080 = { _3573,
                     _2780 };
    assign _3078 = { _3573,
                     _2840 };
    assign _3081 = _3078 + _3080;
    assign _3084 = _3081 + _3083;
    assign _3087 = _3084 + _3086;
    assign _3090 = _3087 + _3089;
    assign _3092 = _3090 < _3576;
    assign _3093 = _2810 & _3092;
    assign _3548 = ~ _3093;
    assign _3549 = _2810 & _3548;
    assign _3550 = _221 ? _3549 : _2810;
    assign _3551 = _531 ? _2840 : _3550;
    assign _195 = _3551;
    always @(posedge _209) begin
        if (_223)
            _2810 <= _2929;
        else
            _2810 <= _195;
    end
    assign _3099 = { _3573,
                     _2810 };
    assign _3097 = { _3573,
                     _2870 };
    assign _3100 = _3097 + _3099;
    assign _3103 = _3100 + _3102;
    assign _3106 = _3103 + _3105;
    assign _3109 = _3106 + _3108;
    assign _3111 = _3109 < _3576;
    assign _3112 = _2840 & _3111;
    assign _3552 = ~ _3112;
    assign _3553 = _2840 & _3552;
    assign _3554 = _221 ? _3553 : _2840;
    assign _3555 = _531 ? _2870 : _3554;
    assign _196 = _3555;
    always @(posedge _209) begin
        if (_223)
            _2840 <= _2929;
        else
            _2840 <= _196;
    end
    assign _3118 = { _3573,
                     _2840 };
    assign _3116 = { _3573,
                     _2900 };
    assign _3119 = _3116 + _3118;
    assign _3122 = _3119 + _3121;
    assign _3125 = _3122 + _3124;
    assign _3128 = _3125 + _3127;
    assign _3130 = _3128 < _3576;
    assign _3131 = _2870 & _3130;
    assign _3556 = ~ _3131;
    assign _3557 = _2870 & _3556;
    assign _3558 = _221 ? _3557 : _2870;
    assign _3559 = _531 ? _2900 : _3558;
    assign _197 = _3559;
    always @(posedge _209) begin
        if (_223)
            _2870 <= _2929;
        else
            _2870 <= _197;
    end
    assign _3137 = { _3573,
                     _2870 };
    assign _3135 = { _3573,
                     _2930 };
    assign _3138 = _3135 + _3137;
    assign _3141 = _3138 + _3140;
    assign _3144 = _3141 + _3143;
    assign _3147 = _3144 + _3146;
    assign _3149 = _3147 < _3576;
    assign _3150 = _2900 & _3149;
    assign _3560 = ~ _3150;
    assign _3561 = _2900 & _3560;
    assign _3562 = _221 ? _3561 : _2900;
    assign _3563 = _531 ? _2930 : _3562;
    assign _198 = _3563;
    always @(posedge _209) begin
        if (_223)
            _2900 <= _2929;
        else
            _2900 <= _198;
    end
    assign _3156 = { _3573,
                     _2900 };
    assign _3154 = { _3573,
                     _2960 };
    assign _3157 = _3154 + _3156;
    assign _3160 = _3157 + _3159;
    assign _3163 = _3160 + _3162;
    assign _3166 = _3163 + _3165;
    assign _3168 = _3166 < _3576;
    assign _3169 = _2930 & _3168;
    assign _3564 = ~ _3169;
    assign _3565 = _2930 & _3564;
    assign _3566 = _221 ? _3565 : _2930;
    assign _3567 = _531 ? _2960 : _3566;
    assign _199 = _3567;
    always @(posedge _209) begin
        if (_223)
            _2930 <= _2929;
        else
            _2930 <= _199;
    end
    assign _3569 = { _3573,
                     _2930 };
    assign _3572 = _3569 + _3571;
    assign _3575 = _3572 + _3574;
    assign _3577 = _3575 < _3576;
    assign _222 = _220[1:1];
    assign _223 = _207 | _222;
    assign _3582 = _211[0:0];
    assign _3579 = ~ _3578;
    assign _3580 = _2960 & _3579;
    assign _3581 = _221 ? _3580 : _2960;
    assign _3583 = _531 ? _3582 : _3581;
    assign _200 = _3583;
    always @(posedge _209) begin
        if (_223)
            _2960 <= _2929;
        else
            _2960 <= _200;
    end
    assign _3578 = _2960 & _3577;
    assign gnd = 1'b0;
    assign _3584 = _221 ? _3578 : gnd;
    assign _529 = 4'b0001;
    assign _530 = _203 == _529;
    assign _531 = _205 & _530;
    assign _3585 = _531 ? gnd : _3584;
    assign _201 = _3585;
    assign _229 = { _3891,
                    _201 };
    assign _232 = _229 + _231;
    assign _235 = _232 + _234;
    assign _238 = _235 + _237;
    assign _241 = _238 + _240;
    assign _244 = _241 + _243;
    assign _247 = _244 + _246;
    assign _250 = _247 + _249;
    assign _253 = _250 + _252;
    assign _256 = _253 + _255;
    assign _259 = _256 + _258;
    assign _262 = _259 + _261;
    assign _265 = _262 + _264;
    assign _268 = _265 + _267;
    assign _271 = _268 + _270;
    assign _274 = _271 + _273;
    assign _277 = _274 + _276;
    assign _280 = _277 + _279;
    assign _283 = _280 + _282;
    assign _286 = _283 + _285;
    assign _289 = _286 + _288;
    assign _292 = _289 + _291;
    assign _295 = _292 + _294;
    assign _298 = _295 + _297;
    assign _301 = _298 + _300;
    assign _304 = _301 + _303;
    assign _307 = _304 + _306;
    assign _310 = _307 + _309;
    assign _313 = _310 + _312;
    assign _316 = _313 + _315;
    assign _319 = _316 + _318;
    assign _322 = _319 + _321;
    assign _325 = _322 + _324;
    assign _328 = _325 + _327;
    assign _331 = _328 + _330;
    assign _334 = _331 + _333;
    assign _337 = _334 + _336;
    assign _340 = _337 + _339;
    assign _343 = _340 + _342;
    assign _346 = _343 + _345;
    assign _349 = _346 + _348;
    assign _352 = _349 + _351;
    assign _355 = _352 + _354;
    assign _358 = _355 + _357;
    assign _361 = _358 + _360;
    assign _364 = _361 + _363;
    assign _367 = _364 + _366;
    assign _370 = _367 + _369;
    assign _373 = _370 + _372;
    assign _376 = _373 + _375;
    assign _379 = _376 + _378;
    assign _382 = _379 + _381;
    assign _385 = _382 + _384;
    assign _388 = _385 + _387;
    assign _391 = _388 + _390;
    assign _394 = _391 + _393;
    assign _397 = _394 + _396;
    assign _400 = _397 + _399;
    assign _403 = _400 + _402;
    assign _406 = _403 + _405;
    assign _409 = _406 + _408;
    assign _412 = _409 + _411;
    assign _415 = _412 + _414;
    assign _418 = _415 + _417;
    assign _421 = _418 + _420;
    assign _424 = _421 + _423;
    assign _427 = _424 + _426;
    assign _430 = _427 + _429;
    assign _433 = _430 + _432;
    assign _436 = _433 + _435;
    assign _439 = _436 + _438;
    assign _442 = _439 + _441;
    assign _445 = _442 + _444;
    assign _448 = _445 + _447;
    assign _451 = _448 + _450;
    assign _454 = _451 + _453;
    assign _457 = _454 + _456;
    assign _460 = _457 + _459;
    assign _463 = _460 + _462;
    assign _466 = _463 + _465;
    assign _469 = _466 + _468;
    assign _472 = _469 + _471;
    assign _475 = _472 + _474;
    assign _478 = _475 + _477;
    assign _481 = _478 + _480;
    assign _484 = _481 + _483;
    assign _487 = _484 + _486;
    assign _490 = _487 + _489;
    assign _493 = _490 + _492;
    assign _496 = _493 + _495;
    assign _499 = _496 + _498;
    assign _502 = _499 + _501;
    assign _505 = _502 + _504;
    assign _508 = _505 + _507;
    assign _511 = _508 + _510;
    assign _514 = _511 + _513;
    assign _517 = _514 + _516;
    assign _520 = _517 + _519;
    assign _523 = _520 + _522;
    assign _526 = _523 + _525;
    assign _3589 = _526 == _3594;
    assign _221 = _220[0:0];
    assign _3590 = _221 & _3589;
    assign _3587 = 31'b0000000000000000000000000000000;
    assign _3591 = { _3587,
                     _3590 };
    assign _3586 = 32'b00000000000000000000000000000000;
    assign _217 = 4'b0000;
    assign _203 = write_addr;
    assign _218 = _203 == _217;
    assign _205 = write_enable;
    assign _219 = _205 & _218;
    assign _207 = clear;
    assign _209 = clock;
    assign _211 = write_data;
    assign _212 = _211;
    always @(posedge _209) begin
        if (_207)
            _220 <= _3586;
        else
            if (_219)
                _220 <= _212;
    end
    assign _214 = read_addr;
    always @* begin
        case (_214)
        0:
            _3895 <= _220;
        1:
            _3895 <= _3586;
        2:
            _3895 <= _3591;
        3:
            _3895 <= _3593;
        default:
            _3895 <= _3894;
        endcase
    end
    assign read_data = _3895;

endmodule
module aoc_solver_top (
    read_addr,
    write_data,
    write_addr,
    write_enable,
    clear,
    clock,
    read_data
);

    input [3:0] read_addr;
    input [31:0] write_data;
    input [3:0] write_addr;
    input write_enable;
    input clear;
    input clock;
    output [31:0] read_data;

    wire [3:0] _2;
    wire [31:0] _4;
    wire [3:0] _6;
    wire _8;
    wire _10;
    wire _12;
    wire [31:0] _15;
    wire [31:0] _13;
    assign _2 = read_addr;
    assign _4 = write_data;
    assign _6 = write_addr;
    assign _8 = write_enable;
    assign _10 = clear;
    assign _12 = clock;
    aoc_solver
        aoc_solver
        ( .clock(_12),
          .clear(_10),
          .write_enable(_8),
          .write_addr(_6),
          .write_data(_4),
          .read_addr(_2),
          .read_data(_15[31:0]) );
    assign _13 = _15;
    assign read_data = _13;

endmodule

