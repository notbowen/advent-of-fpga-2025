module aoc_solver (
    clear,
    clock,
    load_data,
    load,
    start,
    finished,
    total_removed,
    current_active
);

    input clear;
    input clock;
    input load_data;
    input load;
    input start;
    output finished;
    output [15:0] total_removed;
    output [15:0] current_active;

    wire [14:0] _709;
    wire [15:0] _712;
    wire [15:0] _707;
    wire [15:0] _702;
    wire [15:0] _697;
    wire [15:0] _692;
    wire [15:0] _687;
    wire [15:0] _682;
    wire [15:0] _677;
    wire [15:0] _672;
    wire [15:0] _667;
    wire [15:0] _662;
    wire [15:0] _657;
    wire [15:0] _652;
    wire [15:0] _647;
    wire [15:0] _642;
    wire [15:0] _637;
    wire [15:0] _632;
    wire [15:0] _627;
    wire [15:0] _622;
    wire [15:0] _617;
    wire [15:0] _612;
    wire [15:0] _607;
    wire [15:0] _602;
    wire [15:0] _597;
    wire [15:0] _592;
    wire [15:0] _587;
    wire [15:0] _582;
    wire [15:0] _577;
    wire [15:0] _572;
    wire [15:0] _567;
    wire [15:0] _562;
    wire [15:0] _557;
    wire [15:0] _552;
    wire [15:0] _547;
    wire [15:0] _542;
    wire [15:0] _537;
    wire [15:0] _532;
    wire [15:0] _527;
    wire [15:0] _522;
    wire [15:0] _517;
    wire [15:0] _512;
    wire [15:0] _507;
    wire [15:0] _502;
    wire [15:0] _497;
    wire [15:0] _492;
    wire [15:0] _487;
    wire [15:0] _482;
    wire [15:0] _477;
    wire [15:0] _472;
    wire [15:0] _467;
    wire [15:0] _462;
    wire [15:0] _457;
    wire [15:0] _452;
    wire [15:0] _447;
    wire [15:0] _442;
    wire [15:0] _437;
    wire [15:0] _432;
    wire [15:0] _427;
    wire [15:0] _422;
    wire [15:0] _417;
    wire [15:0] _412;
    wire [15:0] _407;
    wire [15:0] _402;
    wire [15:0] _397;
    wire [15:0] _392;
    wire [15:0] _387;
    wire [15:0] _382;
    wire [15:0] _377;
    wire [15:0] _372;
    wire [15:0] _367;
    wire [15:0] _362;
    wire [15:0] _357;
    wire [15:0] _352;
    wire [15:0] _347;
    wire [15:0] _342;
    wire [15:0] _337;
    wire [15:0] _332;
    wire [15:0] _327;
    wire [15:0] _322;
    wire [15:0] _317;
    wire [15:0] _312;
    wire [15:0] _307;
    wire [15:0] _302;
    wire [15:0] _297;
    wire [15:0] _292;
    wire [15:0] _287;
    wire [15:0] _282;
    wire [15:0] _277;
    wire [15:0] _272;
    wire [15:0] _267;
    wire [15:0] _262;
    wire [15:0] _257;
    wire [15:0] _252;
    wire [15:0] _247;
    wire [15:0] _242;
    wire [15:0] _237;
    wire [15:0] _232;
    wire [15:0] _227;
    wire [15:0] _222;
    wire [15:0] _218;
    wire [15:0] _223;
    wire [15:0] _228;
    wire [15:0] _233;
    wire [15:0] _238;
    wire [15:0] _243;
    wire [15:0] _248;
    wire [15:0] _253;
    wire [15:0] _258;
    wire [15:0] _263;
    wire [15:0] _268;
    wire [15:0] _273;
    wire [15:0] _278;
    wire [15:0] _283;
    wire [15:0] _288;
    wire [15:0] _293;
    wire [15:0] _298;
    wire [15:0] _303;
    wire [15:0] _308;
    wire [15:0] _313;
    wire [15:0] _318;
    wire [15:0] _323;
    wire [15:0] _328;
    wire [15:0] _333;
    wire [15:0] _338;
    wire [15:0] _343;
    wire [15:0] _348;
    wire [15:0] _353;
    wire [15:0] _358;
    wire [15:0] _363;
    wire [15:0] _368;
    wire [15:0] _373;
    wire [15:0] _378;
    wire [15:0] _383;
    wire [15:0] _388;
    wire [15:0] _393;
    wire [15:0] _398;
    wire [15:0] _403;
    wire [15:0] _408;
    wire [15:0] _413;
    wire [15:0] _418;
    wire [15:0] _423;
    wire [15:0] _428;
    wire [15:0] _433;
    wire [15:0] _438;
    wire [15:0] _443;
    wire [15:0] _448;
    wire [15:0] _453;
    wire [15:0] _458;
    wire [15:0] _463;
    wire [15:0] _468;
    wire [15:0] _473;
    wire [15:0] _478;
    wire [15:0] _483;
    wire [15:0] _488;
    wire [15:0] _493;
    wire [15:0] _498;
    wire [15:0] _503;
    wire [15:0] _508;
    wire [15:0] _513;
    wire [15:0] _518;
    wire [15:0] _523;
    wire [15:0] _528;
    wire [15:0] _533;
    wire [15:0] _538;
    wire [15:0] _543;
    wire [15:0] _548;
    wire [15:0] _553;
    wire [15:0] _558;
    wire [15:0] _563;
    wire [15:0] _568;
    wire [15:0] _573;
    wire [15:0] _578;
    wire [15:0] _583;
    wire [15:0] _588;
    wire [15:0] _593;
    wire [15:0] _598;
    wire [15:0] _603;
    wire [15:0] _608;
    wire [15:0] _613;
    wire [15:0] _618;
    wire [15:0] _623;
    wire [15:0] _628;
    wire [15:0] _633;
    wire [15:0] _638;
    wire [15:0] _643;
    wire [15:0] _648;
    wire [15:0] _653;
    wire [15:0] _658;
    wire [15:0] _663;
    wire [15:0] _668;
    wire [15:0] _673;
    wire [15:0] _678;
    wire [15:0] _683;
    wire [15:0] _688;
    wire [15:0] _693;
    wire [15:0] _698;
    wire [15:0] _703;
    wire [15:0] _708;
    wire [15:0] _713;
    wire [15:0] _714;
    wire [15:0] _1017;
    wire [15:0] _717;
    wire [15:0] _1018;
    wire [15:0] _2;
    reg [15:0] _715;
    wire _1031;
    wire _1032;
    wire _4;
    wire [15:0] _1015;
    wire _1050;
    wire _1051;
    wire _5;
    wire [15:0] _1012;
    wire _1069;
    wire _1070;
    wire _6;
    wire [15:0] _1009;
    wire _1088;
    wire _1089;
    wire _7;
    wire [15:0] _1006;
    wire _1107;
    wire _1108;
    wire _8;
    wire [15:0] _1003;
    wire _1126;
    wire _1127;
    wire _9;
    wire [15:0] _1000;
    wire _1145;
    wire _1146;
    wire _10;
    wire [15:0] _997;
    wire _1164;
    wire _1165;
    wire _11;
    wire [15:0] _994;
    wire _1183;
    wire _1184;
    wire _12;
    wire [15:0] _991;
    wire _1196;
    wire _1197;
    wire _13;
    wire [15:0] _988;
    wire _1215;
    wire _1216;
    wire _14;
    wire [15:0] _985;
    wire _1243;
    wire _1244;
    wire _15;
    wire [15:0] _982;
    wire _1271;
    wire _1272;
    wire _16;
    wire [15:0] _979;
    wire _1299;
    wire _1300;
    wire _17;
    wire [15:0] _976;
    wire _1327;
    wire _1328;
    wire _18;
    wire [15:0] _973;
    wire _1355;
    wire _1356;
    wire _19;
    wire [15:0] _970;
    wire _1383;
    wire _1384;
    wire _20;
    wire [15:0] _967;
    wire _1411;
    wire _1412;
    wire _21;
    wire [15:0] _964;
    wire _1439;
    wire _1440;
    wire _22;
    wire [15:0] _961;
    wire _1458;
    wire _1459;
    wire _23;
    wire [15:0] _958;
    wire _1477;
    wire _1478;
    wire _24;
    wire [15:0] _955;
    wire _1505;
    wire _1506;
    wire _25;
    wire [15:0] _952;
    wire _1533;
    wire _1534;
    wire _26;
    wire [15:0] _949;
    wire _1561;
    wire _1562;
    wire _27;
    wire [15:0] _946;
    wire _1589;
    wire _1590;
    wire _28;
    wire [15:0] _943;
    wire _1617;
    wire _1618;
    wire _29;
    wire [15:0] _940;
    wire _1645;
    wire _1646;
    wire _30;
    wire [15:0] _937;
    wire _1673;
    wire _1674;
    wire _31;
    wire [15:0] _934;
    wire _1701;
    wire _1702;
    wire _32;
    wire [15:0] _931;
    wire _1720;
    wire _1721;
    wire _33;
    wire [15:0] _928;
    wire _1739;
    wire _1740;
    wire _34;
    wire [15:0] _925;
    wire _1767;
    wire _1768;
    wire _35;
    wire [15:0] _922;
    wire _1795;
    wire _1796;
    wire _36;
    wire [15:0] _919;
    wire _1823;
    wire _1824;
    wire _37;
    wire [15:0] _916;
    wire _1851;
    wire _1852;
    wire _38;
    wire [15:0] _913;
    wire _1879;
    wire _1880;
    wire _39;
    wire [15:0] _910;
    wire _1907;
    wire _1908;
    wire _40;
    wire [15:0] _907;
    wire _1935;
    wire _1936;
    wire _41;
    wire [15:0] _904;
    wire _1963;
    wire _1964;
    wire _42;
    wire [15:0] _901;
    wire _1982;
    wire _1983;
    wire _43;
    wire [15:0] _898;
    wire _2001;
    wire _2002;
    wire _44;
    wire [15:0] _895;
    wire _2029;
    wire _2030;
    wire _45;
    wire [15:0] _892;
    wire _2057;
    wire _2058;
    wire _46;
    wire [15:0] _889;
    wire _2085;
    wire _2086;
    wire _47;
    wire [15:0] _886;
    wire _2113;
    wire _2114;
    wire _48;
    wire [15:0] _883;
    wire _2141;
    wire _2142;
    wire _49;
    wire [15:0] _880;
    wire _2169;
    wire _2170;
    wire _50;
    wire [15:0] _877;
    wire _2197;
    wire _2198;
    wire _51;
    wire [15:0] _874;
    wire _2225;
    wire _2226;
    wire _52;
    wire [15:0] _871;
    wire _2244;
    wire _2245;
    wire _53;
    wire [15:0] _868;
    wire _2263;
    wire _2264;
    wire _54;
    wire [15:0] _865;
    wire _2291;
    wire _2292;
    wire _55;
    wire [15:0] _862;
    wire _2319;
    wire _2320;
    wire _56;
    wire [15:0] _859;
    wire _2347;
    wire _2348;
    wire _57;
    wire [15:0] _856;
    wire _2375;
    wire _2376;
    wire _58;
    wire [15:0] _853;
    wire _2403;
    wire _2404;
    wire _59;
    wire [15:0] _850;
    wire _2431;
    wire _2432;
    wire _60;
    wire [15:0] _847;
    wire _2459;
    wire _2460;
    wire _61;
    wire [15:0] _844;
    wire _2487;
    wire _2488;
    wire _62;
    wire [15:0] _841;
    wire _2506;
    wire _2507;
    wire _63;
    wire [15:0] _838;
    wire _2525;
    wire _2526;
    wire _64;
    wire [15:0] _835;
    wire _2553;
    wire _2554;
    wire _65;
    wire [15:0] _832;
    wire _2581;
    wire _2582;
    wire _66;
    wire [15:0] _829;
    wire _2609;
    wire _2610;
    wire _67;
    wire [15:0] _826;
    wire _2637;
    wire _2638;
    wire _68;
    wire [15:0] _823;
    wire _2665;
    wire _2666;
    wire _69;
    wire [15:0] _820;
    wire _2693;
    wire _2694;
    wire _70;
    wire [15:0] _817;
    wire _2721;
    wire _2722;
    wire _71;
    wire [15:0] _814;
    wire _2749;
    wire _2750;
    wire _72;
    wire [15:0] _811;
    wire _2768;
    wire _2769;
    wire _73;
    wire [15:0] _808;
    wire _2787;
    wire _2788;
    wire _74;
    wire [15:0] _805;
    wire _2815;
    wire _2816;
    wire _75;
    wire [15:0] _802;
    wire _2843;
    wire _2844;
    wire _76;
    wire [15:0] _799;
    wire _2871;
    wire _2872;
    wire _77;
    wire [15:0] _796;
    wire _2899;
    wire _2900;
    wire _78;
    wire [15:0] _793;
    wire _2927;
    wire _2928;
    wire _79;
    wire [15:0] _790;
    wire _2955;
    wire _2956;
    wire _80;
    wire [15:0] _787;
    wire _2983;
    wire _2984;
    wire _81;
    wire [15:0] _784;
    wire _3011;
    wire _3012;
    wire _82;
    wire [15:0] _781;
    wire _3030;
    wire _3031;
    wire _83;
    wire [15:0] _778;
    wire _3049;
    wire _3050;
    wire _84;
    wire [15:0] _775;
    wire _3077;
    wire _3078;
    wire _85;
    wire [15:0] _772;
    wire _3105;
    wire _3106;
    wire _86;
    wire [15:0] _769;
    wire _3133;
    wire _3134;
    wire _87;
    wire [15:0] _766;
    wire _3161;
    wire _3162;
    wire _88;
    wire [15:0] _763;
    wire _3189;
    wire _3190;
    wire _89;
    wire [15:0] _760;
    wire _3217;
    wire _3218;
    wire _90;
    wire [15:0] _757;
    wire _3245;
    wire _3246;
    wire _91;
    wire [15:0] _754;
    wire _3273;
    wire _3274;
    wire _92;
    wire [15:0] _751;
    wire _3292;
    wire _3293;
    wire _93;
    wire [15:0] _748;
    wire _3305;
    wire _3306;
    wire _94;
    wire [15:0] _745;
    wire _3324;
    wire _3325;
    wire _95;
    wire [15:0] _742;
    wire _3343;
    wire _3344;
    wire _96;
    wire [15:0] _739;
    wire _3362;
    wire _3363;
    wire _97;
    wire [15:0] _736;
    wire _3381;
    wire _3382;
    wire _98;
    wire [15:0] _733;
    wire _3400;
    wire _3401;
    wire _99;
    wire [15:0] _730;
    wire _3419;
    wire _3420;
    wire _100;
    wire [15:0] _727;
    wire _3438;
    wire _3439;
    wire _101;
    wire [15:0] _724;
    wire _3457;
    wire _3458;
    wire _102;
    wire [15:0] _721;
    wire [3:0] _3863;
    wire [2:0] _3860;
    wire [3:0] _3861;
    wire [3:0] _3858;
    wire _220;
    wire [3:0] _3452;
    wire [3:0] _3449;
    wire [3:0] _3446;
    wire [3:0] _3433;
    wire [3:0] _3430;
    wire [3:0] _3427;
    wire [3:0] _3414;
    wire [3:0] _3411;
    wire [3:0] _3408;
    wire [3:0] _3395;
    wire [3:0] _3392;
    wire [3:0] _3389;
    wire [3:0] _3376;
    wire [3:0] _3373;
    wire [3:0] _3370;
    wire [3:0] _3357;
    wire [3:0] _3354;
    wire [3:0] _3351;
    wire [3:0] _3338;
    wire [3:0] _3335;
    wire [3:0] _3332;
    wire [3:0] _3319;
    wire [3:0] _3316;
    wire [3:0] _3313;
    wire [3:0] _3300;
    wire [3:0] _3072;
    wire [3:0] _3069;
    wire [3:0] _3066;
    wire [3:0] _3063;
    wire [3:0] _3100;
    wire [3:0] _3097;
    wire [3:0] _3094;
    wire [3:0] _3091;
    wire [3:0] _3128;
    wire [3:0] _3125;
    wire [3:0] _3122;
    wire [3:0] _3119;
    wire [3:0] _3156;
    wire [3:0] _3153;
    wire [3:0] _3150;
    wire [3:0] _3147;
    wire [3:0] _3184;
    wire [3:0] _3181;
    wire [3:0] _3178;
    wire [3:0] _3175;
    wire [3:0] _3212;
    wire [3:0] _3209;
    wire [3:0] _3206;
    wire [3:0] _3203;
    wire [3:0] _3240;
    wire [3:0] _3237;
    wire [3:0] _3234;
    wire [3:0] _3231;
    wire [3:0] _3268;
    wire [3:0] _3265;
    wire [3:0] _3262;
    wire [3:0] _3259;
    wire [3:0] _3287;
    wire [3:0] _3025;
    wire [3:0] _3022;
    wire [3:0] _3006;
    wire [3:0] _3003;
    wire [3:0] _3000;
    wire [3:0] _2978;
    wire [3:0] _2975;
    wire [3:0] _2972;
    wire [3:0] _2950;
    wire [3:0] _2947;
    wire [3:0] _2944;
    wire [3:0] _2922;
    wire [3:0] _2919;
    wire [3:0] _2916;
    wire [3:0] _2894;
    wire [3:0] _2891;
    wire [3:0] _2888;
    wire [3:0] _2866;
    wire [3:0] _2863;
    wire [3:0] _2860;
    wire [3:0] _2838;
    wire [3:0] _2835;
    wire [3:0] _2832;
    wire [3:0] _2810;
    wire [3:0] _2807;
    wire [3:0] _2804;
    wire [3:0] _2801;
    wire [3:0] _2798;
    wire [3:0] _2782;
    wire [3:0] _2548;
    wire [3:0] _2545;
    wire [3:0] _2542;
    wire [3:0] _2539;
    wire [3:0] _2576;
    wire [3:0] _2573;
    wire [3:0] _2570;
    wire [3:0] _2567;
    wire [3:0] _2604;
    wire [3:0] _2601;
    wire [3:0] _2598;
    wire [3:0] _2595;
    wire [3:0] _2632;
    wire [3:0] _2629;
    wire [3:0] _2626;
    wire [3:0] _2623;
    wire [3:0] _2660;
    wire [3:0] _2657;
    wire [3:0] _2654;
    wire [3:0] _2651;
    wire [3:0] _2688;
    wire [3:0] _2685;
    wire [3:0] _2682;
    wire [3:0] _2679;
    wire [3:0] _2716;
    wire [3:0] _2713;
    wire [3:0] _2710;
    wire [3:0] _2707;
    wire [3:0] _2744;
    wire [3:0] _2741;
    wire [3:0] _2738;
    wire [3:0] _2735;
    wire [3:0] _2763;
    wire [3:0] _2501;
    wire [3:0] _2498;
    wire [3:0] _2482;
    wire [3:0] _2479;
    wire [3:0] _2476;
    wire [3:0] _2454;
    wire [3:0] _2451;
    wire [3:0] _2448;
    wire [3:0] _2426;
    wire [3:0] _2423;
    wire [3:0] _2420;
    wire [3:0] _2398;
    wire [3:0] _2395;
    wire [3:0] _2392;
    wire [3:0] _2370;
    wire [3:0] _2367;
    wire [3:0] _2364;
    wire [3:0] _2342;
    wire [3:0] _2339;
    wire [3:0] _2336;
    wire [3:0] _2314;
    wire [3:0] _2311;
    wire [3:0] _2308;
    wire [3:0] _2286;
    wire [3:0] _2283;
    wire [3:0] _2280;
    wire [3:0] _2277;
    wire [3:0] _2274;
    wire [3:0] _2258;
    wire [3:0] _2024;
    wire [3:0] _2021;
    wire [3:0] _2018;
    wire [3:0] _2015;
    wire [3:0] _2052;
    wire [3:0] _2049;
    wire [3:0] _2046;
    wire [3:0] _2043;
    wire [3:0] _2080;
    wire [3:0] _2077;
    wire [3:0] _2074;
    wire [3:0] _2071;
    wire [3:0] _2108;
    wire [3:0] _2105;
    wire [3:0] _2102;
    wire [3:0] _2099;
    wire [3:0] _2136;
    wire [3:0] _2133;
    wire [3:0] _2130;
    wire [3:0] _2127;
    wire [3:0] _2164;
    wire [3:0] _2161;
    wire [3:0] _2158;
    wire [3:0] _2155;
    wire [3:0] _2192;
    wire [3:0] _2189;
    wire [3:0] _2186;
    wire [3:0] _2183;
    wire [3:0] _2220;
    wire [3:0] _2217;
    wire [3:0] _2214;
    wire [3:0] _2211;
    wire [3:0] _2239;
    wire [3:0] _1977;
    wire [3:0] _1974;
    wire [3:0] _1958;
    wire [3:0] _1955;
    wire [3:0] _1952;
    wire [3:0] _1930;
    wire [3:0] _1927;
    wire [3:0] _1924;
    wire [3:0] _1902;
    wire [3:0] _1899;
    wire [3:0] _1896;
    wire [3:0] _1874;
    wire [3:0] _1871;
    wire [3:0] _1868;
    wire [3:0] _1846;
    wire [3:0] _1843;
    wire [3:0] _1840;
    wire [3:0] _1818;
    wire [3:0] _1815;
    wire [3:0] _1812;
    wire [3:0] _1790;
    wire [3:0] _1787;
    wire [3:0] _1784;
    wire [3:0] _1762;
    wire [3:0] _1759;
    wire [3:0] _1756;
    wire [3:0] _1753;
    wire [3:0] _1750;
    wire [3:0] _1734;
    wire [3:0] _1500;
    wire [3:0] _1497;
    wire [3:0] _1494;
    wire [3:0] _1491;
    wire [3:0] _1528;
    wire [3:0] _1525;
    wire [3:0] _1522;
    wire [3:0] _1519;
    wire [3:0] _1556;
    wire [3:0] _1553;
    wire [3:0] _1550;
    wire [3:0] _1547;
    wire [3:0] _1584;
    wire [3:0] _1581;
    wire [3:0] _1578;
    wire [3:0] _1575;
    wire [3:0] _1612;
    wire [3:0] _1609;
    wire [3:0] _1606;
    wire [3:0] _1603;
    wire [3:0] _1640;
    wire [3:0] _1637;
    wire [3:0] _1634;
    wire [3:0] _1631;
    wire [3:0] _1668;
    wire [3:0] _1665;
    wire [3:0] _1662;
    wire [3:0] _1659;
    wire [3:0] _1696;
    wire [3:0] _1693;
    wire [3:0] _1690;
    wire [3:0] _1687;
    wire [3:0] _1715;
    wire [3:0] _1453;
    wire [3:0] _1450;
    wire [3:0] _1434;
    wire [3:0] _1431;
    wire [3:0] _1428;
    wire [3:0] _1406;
    wire [3:0] _1403;
    wire [3:0] _1400;
    wire [3:0] _1378;
    wire [3:0] _1375;
    wire [3:0] _1372;
    wire [3:0] _1350;
    wire [3:0] _1347;
    wire [3:0] _1344;
    wire [3:0] _1322;
    wire [3:0] _1319;
    wire [3:0] _1316;
    wire [3:0] _1294;
    wire [3:0] _1291;
    wire [3:0] _1288;
    wire [3:0] _1266;
    wire [3:0] _1263;
    wire [3:0] _1260;
    wire [3:0] _1238;
    wire [3:0] _1235;
    wire [3:0] _1232;
    wire [3:0] _1229;
    wire [3:0] _1226;
    wire [3:0] _1210;
    wire [3:0] _1026;
    wire [3:0] _1023;
    wire [3:0] _1021;
    wire [3:0] _1024;
    wire [3:0] _1027;
    wire _1029;
    wire _1030;
    wire _3459;
    wire _3460;
    wire _3461;
    wire _3462;
    wire _103;
    reg _711;
    wire [3:0] _1045;
    wire [3:0] _1064;
    wire [3:0] _1083;
    wire [3:0] _1102;
    wire [3:0] _1121;
    wire [3:0] _1140;
    wire [3:0] _1159;
    wire [3:0] _1178;
    wire [3:0] _1191;
    wire [3:0] _1188;
    wire [3:0] _1186;
    wire [3:0] _1189;
    wire [3:0] _1192;
    wire _1194;
    wire _1195;
    wire _3463;
    wire _3464;
    wire _3465;
    wire _3466;
    wire _104;
    reg _666;
    wire [3:0] _1175;
    wire [3:0] _1172;
    wire [3:0] _1169;
    wire [3:0] _1167;
    wire [3:0] _1170;
    wire [3:0] _1173;
    wire [3:0] _1176;
    wire [3:0] _1179;
    wire _1181;
    wire _1182;
    wire _3467;
    wire _3468;
    wire _3469;
    wire _3470;
    wire _105;
    reg _671;
    wire [3:0] _1156;
    wire [3:0] _1153;
    wire [3:0] _1150;
    wire [3:0] _1148;
    wire [3:0] _1151;
    wire [3:0] _1154;
    wire [3:0] _1157;
    wire [3:0] _1160;
    wire _1162;
    wire _1163;
    wire _3471;
    wire _3472;
    wire _3473;
    wire _3474;
    wire _106;
    reg _676;
    wire [3:0] _1137;
    wire [3:0] _1134;
    wire [3:0] _1131;
    wire [3:0] _1129;
    wire [3:0] _1132;
    wire [3:0] _1135;
    wire [3:0] _1138;
    wire [3:0] _1141;
    wire _1143;
    wire _1144;
    wire _3475;
    wire _3476;
    wire _3477;
    wire _3478;
    wire _107;
    reg _681;
    wire [3:0] _1118;
    wire [3:0] _1115;
    wire [3:0] _1112;
    wire [3:0] _1110;
    wire [3:0] _1113;
    wire [3:0] _1116;
    wire [3:0] _1119;
    wire [3:0] _1122;
    wire _1124;
    wire _1125;
    wire _3479;
    wire _3480;
    wire _3481;
    wire _3482;
    wire _108;
    reg _686;
    wire [3:0] _1099;
    wire [3:0] _1096;
    wire [3:0] _1093;
    wire [3:0] _1091;
    wire [3:0] _1094;
    wire [3:0] _1097;
    wire [3:0] _1100;
    wire [3:0] _1103;
    wire _1105;
    wire _1106;
    wire _3483;
    wire _3484;
    wire _3485;
    wire _3486;
    wire _109;
    reg _691;
    wire [3:0] _1080;
    wire [3:0] _1077;
    wire [3:0] _1074;
    wire [3:0] _1072;
    wire [3:0] _1075;
    wire [3:0] _1078;
    wire [3:0] _1081;
    wire [3:0] _1084;
    wire _1086;
    wire _1087;
    wire _3487;
    wire _3488;
    wire _3489;
    wire _3490;
    wire _110;
    reg _696;
    wire [3:0] _1061;
    wire [3:0] _1058;
    wire [3:0] _1055;
    wire [3:0] _1053;
    wire [3:0] _1056;
    wire [3:0] _1059;
    wire [3:0] _1062;
    wire [3:0] _1065;
    wire _1067;
    wire _1068;
    wire _3491;
    wire _3492;
    wire _3493;
    wire _3494;
    wire _111;
    reg _701;
    wire [3:0] _1042;
    wire [3:0] _1039;
    wire [3:0] _1036;
    wire [3:0] _1034;
    wire [3:0] _1037;
    wire [3:0] _1040;
    wire [3:0] _1043;
    wire [3:0] _1046;
    wire _1048;
    wire _1049;
    wire _3495;
    wire _3496;
    wire _3497;
    wire _3498;
    wire _112;
    reg _706;
    wire [3:0] _1207;
    wire [3:0] _1204;
    wire [3:0] _1201;
    wire [3:0] _1199;
    wire [3:0] _1202;
    wire [3:0] _1205;
    wire [3:0] _1208;
    wire [3:0] _1211;
    wire _1213;
    wire _1214;
    wire _3499;
    wire _3500;
    wire _3501;
    wire _3502;
    wire _113;
    reg _661;
    wire [3:0] _1472;
    wire [3:0] _1469;
    wire [3:0] _1466;
    wire [3:0] _1463;
    wire [3:0] _1461;
    wire [3:0] _1464;
    wire [3:0] _1467;
    wire [3:0] _1470;
    wire [3:0] _1473;
    wire _1475;
    wire _1476;
    wire _3503;
    wire _3504;
    wire _3505;
    wire _3506;
    wire _114;
    reg _611;
    wire [3:0] _1223;
    wire [3:0] _1220;
    wire [3:0] _1218;
    wire [3:0] _1221;
    wire [3:0] _1224;
    wire [3:0] _1227;
    wire [3:0] _1230;
    wire [3:0] _1233;
    wire [3:0] _1236;
    wire [3:0] _1239;
    wire _1241;
    wire _1242;
    wire _3507;
    wire _3508;
    wire _3509;
    wire _3510;
    wire _115;
    reg _656;
    wire [3:0] _1257;
    wire [3:0] _1254;
    wire [3:0] _1251;
    wire [3:0] _1248;
    wire [3:0] _1246;
    wire [3:0] _1249;
    wire [3:0] _1252;
    wire [3:0] _1255;
    wire [3:0] _1258;
    wire [3:0] _1261;
    wire [3:0] _1264;
    wire [3:0] _1267;
    wire _1269;
    wire _1270;
    wire _3511;
    wire _3512;
    wire _3513;
    wire _3514;
    wire _116;
    reg _651;
    wire [3:0] _1285;
    wire [3:0] _1282;
    wire [3:0] _1279;
    wire [3:0] _1276;
    wire [3:0] _1274;
    wire [3:0] _1277;
    wire [3:0] _1280;
    wire [3:0] _1283;
    wire [3:0] _1286;
    wire [3:0] _1289;
    wire [3:0] _1292;
    wire [3:0] _1295;
    wire _1297;
    wire _1298;
    wire _3515;
    wire _3516;
    wire _3517;
    wire _3518;
    wire _117;
    reg _646;
    wire [3:0] _1313;
    wire [3:0] _1310;
    wire [3:0] _1307;
    wire [3:0] _1304;
    wire [3:0] _1302;
    wire [3:0] _1305;
    wire [3:0] _1308;
    wire [3:0] _1311;
    wire [3:0] _1314;
    wire [3:0] _1317;
    wire [3:0] _1320;
    wire [3:0] _1323;
    wire _1325;
    wire _1326;
    wire _3519;
    wire _3520;
    wire _3521;
    wire _3522;
    wire _118;
    reg _641;
    wire [3:0] _1341;
    wire [3:0] _1338;
    wire [3:0] _1335;
    wire [3:0] _1332;
    wire [3:0] _1330;
    wire [3:0] _1333;
    wire [3:0] _1336;
    wire [3:0] _1339;
    wire [3:0] _1342;
    wire [3:0] _1345;
    wire [3:0] _1348;
    wire [3:0] _1351;
    wire _1353;
    wire _1354;
    wire _3523;
    wire _3524;
    wire _3525;
    wire _3526;
    wire _119;
    reg _636;
    wire [3:0] _1369;
    wire [3:0] _1366;
    wire [3:0] _1363;
    wire [3:0] _1360;
    wire [3:0] _1358;
    wire [3:0] _1361;
    wire [3:0] _1364;
    wire [3:0] _1367;
    wire [3:0] _1370;
    wire [3:0] _1373;
    wire [3:0] _1376;
    wire [3:0] _1379;
    wire _1381;
    wire _1382;
    wire _3527;
    wire _3528;
    wire _3529;
    wire _3530;
    wire _120;
    reg _631;
    wire [3:0] _1397;
    wire [3:0] _1394;
    wire [3:0] _1391;
    wire [3:0] _1388;
    wire [3:0] _1386;
    wire [3:0] _1389;
    wire [3:0] _1392;
    wire [3:0] _1395;
    wire [3:0] _1398;
    wire [3:0] _1401;
    wire [3:0] _1404;
    wire [3:0] _1407;
    wire _1409;
    wire _1410;
    wire _3531;
    wire _3532;
    wire _3533;
    wire _3534;
    wire _121;
    reg _626;
    wire [3:0] _1425;
    wire [3:0] _1422;
    wire [3:0] _1419;
    wire [3:0] _1416;
    wire [3:0] _1414;
    wire [3:0] _1417;
    wire [3:0] _1420;
    wire [3:0] _1423;
    wire [3:0] _1426;
    wire [3:0] _1429;
    wire [3:0] _1432;
    wire [3:0] _1435;
    wire _1437;
    wire _1438;
    wire _3535;
    wire _3536;
    wire _3537;
    wire _3538;
    wire _122;
    reg _621;
    wire [3:0] _1447;
    wire [3:0] _1444;
    wire [3:0] _1442;
    wire [3:0] _1445;
    wire [3:0] _1448;
    wire [3:0] _1451;
    wire [3:0] _1454;
    wire _1456;
    wire _1457;
    wire _3539;
    wire _3540;
    wire _3541;
    wire _3542;
    wire _123;
    reg _616;
    wire [3:0] _1712;
    wire [3:0] _1709;
    wire [3:0] _1706;
    wire [3:0] _1704;
    wire [3:0] _1707;
    wire [3:0] _1710;
    wire [3:0] _1713;
    wire [3:0] _1716;
    wire _1718;
    wire _1719;
    wire _3543;
    wire _3544;
    wire _3545;
    wire _3546;
    wire _124;
    reg _566;
    wire [3:0] _1684;
    wire [3:0] _1681;
    wire [3:0] _1678;
    wire [3:0] _1676;
    wire [3:0] _1679;
    wire [3:0] _1682;
    wire [3:0] _1685;
    wire [3:0] _1688;
    wire [3:0] _1691;
    wire [3:0] _1694;
    wire [3:0] _1697;
    wire _1699;
    wire _1700;
    wire _3547;
    wire _3548;
    wire _3549;
    wire _3550;
    wire _125;
    reg _571;
    wire [3:0] _1656;
    wire [3:0] _1653;
    wire [3:0] _1650;
    wire [3:0] _1648;
    wire [3:0] _1651;
    wire [3:0] _1654;
    wire [3:0] _1657;
    wire [3:0] _1660;
    wire [3:0] _1663;
    wire [3:0] _1666;
    wire [3:0] _1669;
    wire _1671;
    wire _1672;
    wire _3551;
    wire _3552;
    wire _3553;
    wire _3554;
    wire _126;
    reg _576;
    wire [3:0] _1628;
    wire [3:0] _1625;
    wire [3:0] _1622;
    wire [3:0] _1620;
    wire [3:0] _1623;
    wire [3:0] _1626;
    wire [3:0] _1629;
    wire [3:0] _1632;
    wire [3:0] _1635;
    wire [3:0] _1638;
    wire [3:0] _1641;
    wire _1643;
    wire _1644;
    wire _3555;
    wire _3556;
    wire _3557;
    wire _3558;
    wire _127;
    reg _581;
    wire [3:0] _1600;
    wire [3:0] _1597;
    wire [3:0] _1594;
    wire [3:0] _1592;
    wire [3:0] _1595;
    wire [3:0] _1598;
    wire [3:0] _1601;
    wire [3:0] _1604;
    wire [3:0] _1607;
    wire [3:0] _1610;
    wire [3:0] _1613;
    wire _1615;
    wire _1616;
    wire _3559;
    wire _3560;
    wire _3561;
    wire _3562;
    wire _128;
    reg _586;
    wire [3:0] _1572;
    wire [3:0] _1569;
    wire [3:0] _1566;
    wire [3:0] _1564;
    wire [3:0] _1567;
    wire [3:0] _1570;
    wire [3:0] _1573;
    wire [3:0] _1576;
    wire [3:0] _1579;
    wire [3:0] _1582;
    wire [3:0] _1585;
    wire _1587;
    wire _1588;
    wire _3563;
    wire _3564;
    wire _3565;
    wire _3566;
    wire _129;
    reg _591;
    wire [3:0] _1544;
    wire [3:0] _1541;
    wire [3:0] _1538;
    wire [3:0] _1536;
    wire [3:0] _1539;
    wire [3:0] _1542;
    wire [3:0] _1545;
    wire [3:0] _1548;
    wire [3:0] _1551;
    wire [3:0] _1554;
    wire [3:0] _1557;
    wire _1559;
    wire _1560;
    wire _3567;
    wire _3568;
    wire _3569;
    wire _3570;
    wire _130;
    reg _596;
    wire [3:0] _1516;
    wire [3:0] _1513;
    wire [3:0] _1510;
    wire [3:0] _1508;
    wire [3:0] _1511;
    wire [3:0] _1514;
    wire [3:0] _1517;
    wire [3:0] _1520;
    wire [3:0] _1523;
    wire [3:0] _1526;
    wire [3:0] _1529;
    wire _1531;
    wire _1532;
    wire _3571;
    wire _3572;
    wire _3573;
    wire _3574;
    wire _131;
    reg _601;
    wire [3:0] _1488;
    wire [3:0] _1485;
    wire [3:0] _1482;
    wire [3:0] _1480;
    wire [3:0] _1483;
    wire [3:0] _1486;
    wire [3:0] _1489;
    wire [3:0] _1492;
    wire [3:0] _1495;
    wire [3:0] _1498;
    wire [3:0] _1501;
    wire _1503;
    wire _1504;
    wire _3575;
    wire _3576;
    wire _3577;
    wire _3578;
    wire _132;
    reg _606;
    wire [3:0] _1731;
    wire [3:0] _1728;
    wire [3:0] _1725;
    wire [3:0] _1723;
    wire [3:0] _1726;
    wire [3:0] _1729;
    wire [3:0] _1732;
    wire [3:0] _1735;
    wire _1737;
    wire _1738;
    wire _3579;
    wire _3580;
    wire _3581;
    wire _3582;
    wire _133;
    reg _561;
    wire [3:0] _1996;
    wire [3:0] _1993;
    wire [3:0] _1990;
    wire [3:0] _1987;
    wire [3:0] _1985;
    wire [3:0] _1988;
    wire [3:0] _1991;
    wire [3:0] _1994;
    wire [3:0] _1997;
    wire _1999;
    wire _2000;
    wire _3583;
    wire _3584;
    wire _3585;
    wire _3586;
    wire _134;
    reg _511;
    wire [3:0] _1747;
    wire [3:0] _1744;
    wire [3:0] _1742;
    wire [3:0] _1745;
    wire [3:0] _1748;
    wire [3:0] _1751;
    wire [3:0] _1754;
    wire [3:0] _1757;
    wire [3:0] _1760;
    wire [3:0] _1763;
    wire _1765;
    wire _1766;
    wire _3587;
    wire _3588;
    wire _3589;
    wire _3590;
    wire _135;
    reg _556;
    wire [3:0] _1781;
    wire [3:0] _1778;
    wire [3:0] _1775;
    wire [3:0] _1772;
    wire [3:0] _1770;
    wire [3:0] _1773;
    wire [3:0] _1776;
    wire [3:0] _1779;
    wire [3:0] _1782;
    wire [3:0] _1785;
    wire [3:0] _1788;
    wire [3:0] _1791;
    wire _1793;
    wire _1794;
    wire _3591;
    wire _3592;
    wire _3593;
    wire _3594;
    wire _136;
    reg _551;
    wire [3:0] _1809;
    wire [3:0] _1806;
    wire [3:0] _1803;
    wire [3:0] _1800;
    wire [3:0] _1798;
    wire [3:0] _1801;
    wire [3:0] _1804;
    wire [3:0] _1807;
    wire [3:0] _1810;
    wire [3:0] _1813;
    wire [3:0] _1816;
    wire [3:0] _1819;
    wire _1821;
    wire _1822;
    wire _3595;
    wire _3596;
    wire _3597;
    wire _3598;
    wire _137;
    reg _546;
    wire [3:0] _1837;
    wire [3:0] _1834;
    wire [3:0] _1831;
    wire [3:0] _1828;
    wire [3:0] _1826;
    wire [3:0] _1829;
    wire [3:0] _1832;
    wire [3:0] _1835;
    wire [3:0] _1838;
    wire [3:0] _1841;
    wire [3:0] _1844;
    wire [3:0] _1847;
    wire _1849;
    wire _1850;
    wire _3599;
    wire _3600;
    wire _3601;
    wire _3602;
    wire _138;
    reg _541;
    wire [3:0] _1865;
    wire [3:0] _1862;
    wire [3:0] _1859;
    wire [3:0] _1856;
    wire [3:0] _1854;
    wire [3:0] _1857;
    wire [3:0] _1860;
    wire [3:0] _1863;
    wire [3:0] _1866;
    wire [3:0] _1869;
    wire [3:0] _1872;
    wire [3:0] _1875;
    wire _1877;
    wire _1878;
    wire _3603;
    wire _3604;
    wire _3605;
    wire _3606;
    wire _139;
    reg _536;
    wire [3:0] _1893;
    wire [3:0] _1890;
    wire [3:0] _1887;
    wire [3:0] _1884;
    wire [3:0] _1882;
    wire [3:0] _1885;
    wire [3:0] _1888;
    wire [3:0] _1891;
    wire [3:0] _1894;
    wire [3:0] _1897;
    wire [3:0] _1900;
    wire [3:0] _1903;
    wire _1905;
    wire _1906;
    wire _3607;
    wire _3608;
    wire _3609;
    wire _3610;
    wire _140;
    reg _531;
    wire [3:0] _1921;
    wire [3:0] _1918;
    wire [3:0] _1915;
    wire [3:0] _1912;
    wire [3:0] _1910;
    wire [3:0] _1913;
    wire [3:0] _1916;
    wire [3:0] _1919;
    wire [3:0] _1922;
    wire [3:0] _1925;
    wire [3:0] _1928;
    wire [3:0] _1931;
    wire _1933;
    wire _1934;
    wire _3611;
    wire _3612;
    wire _3613;
    wire _3614;
    wire _141;
    reg _526;
    wire [3:0] _1949;
    wire [3:0] _1946;
    wire [3:0] _1943;
    wire [3:0] _1940;
    wire [3:0] _1938;
    wire [3:0] _1941;
    wire [3:0] _1944;
    wire [3:0] _1947;
    wire [3:0] _1950;
    wire [3:0] _1953;
    wire [3:0] _1956;
    wire [3:0] _1959;
    wire _1961;
    wire _1962;
    wire _3615;
    wire _3616;
    wire _3617;
    wire _3618;
    wire _142;
    reg _521;
    wire [3:0] _1971;
    wire [3:0] _1968;
    wire [3:0] _1966;
    wire [3:0] _1969;
    wire [3:0] _1972;
    wire [3:0] _1975;
    wire [3:0] _1978;
    wire _1980;
    wire _1981;
    wire _3619;
    wire _3620;
    wire _3621;
    wire _3622;
    wire _143;
    reg _516;
    wire [3:0] _2236;
    wire [3:0] _2233;
    wire [3:0] _2230;
    wire [3:0] _2228;
    wire [3:0] _2231;
    wire [3:0] _2234;
    wire [3:0] _2237;
    wire [3:0] _2240;
    wire _2242;
    wire _2243;
    wire _3623;
    wire _3624;
    wire _3625;
    wire _3626;
    wire _144;
    reg _466;
    wire [3:0] _2208;
    wire [3:0] _2205;
    wire [3:0] _2202;
    wire [3:0] _2200;
    wire [3:0] _2203;
    wire [3:0] _2206;
    wire [3:0] _2209;
    wire [3:0] _2212;
    wire [3:0] _2215;
    wire [3:0] _2218;
    wire [3:0] _2221;
    wire _2223;
    wire _2224;
    wire _3627;
    wire _3628;
    wire _3629;
    wire _3630;
    wire _145;
    reg _471;
    wire [3:0] _2180;
    wire [3:0] _2177;
    wire [3:0] _2174;
    wire [3:0] _2172;
    wire [3:0] _2175;
    wire [3:0] _2178;
    wire [3:0] _2181;
    wire [3:0] _2184;
    wire [3:0] _2187;
    wire [3:0] _2190;
    wire [3:0] _2193;
    wire _2195;
    wire _2196;
    wire _3631;
    wire _3632;
    wire _3633;
    wire _3634;
    wire _146;
    reg _476;
    wire [3:0] _2152;
    wire [3:0] _2149;
    wire [3:0] _2146;
    wire [3:0] _2144;
    wire [3:0] _2147;
    wire [3:0] _2150;
    wire [3:0] _2153;
    wire [3:0] _2156;
    wire [3:0] _2159;
    wire [3:0] _2162;
    wire [3:0] _2165;
    wire _2167;
    wire _2168;
    wire _3635;
    wire _3636;
    wire _3637;
    wire _3638;
    wire _147;
    reg _481;
    wire [3:0] _2124;
    wire [3:0] _2121;
    wire [3:0] _2118;
    wire [3:0] _2116;
    wire [3:0] _2119;
    wire [3:0] _2122;
    wire [3:0] _2125;
    wire [3:0] _2128;
    wire [3:0] _2131;
    wire [3:0] _2134;
    wire [3:0] _2137;
    wire _2139;
    wire _2140;
    wire _3639;
    wire _3640;
    wire _3641;
    wire _3642;
    wire _148;
    reg _486;
    wire [3:0] _2096;
    wire [3:0] _2093;
    wire [3:0] _2090;
    wire [3:0] _2088;
    wire [3:0] _2091;
    wire [3:0] _2094;
    wire [3:0] _2097;
    wire [3:0] _2100;
    wire [3:0] _2103;
    wire [3:0] _2106;
    wire [3:0] _2109;
    wire _2111;
    wire _2112;
    wire _3643;
    wire _3644;
    wire _3645;
    wire _3646;
    wire _149;
    reg _491;
    wire [3:0] _2068;
    wire [3:0] _2065;
    wire [3:0] _2062;
    wire [3:0] _2060;
    wire [3:0] _2063;
    wire [3:0] _2066;
    wire [3:0] _2069;
    wire [3:0] _2072;
    wire [3:0] _2075;
    wire [3:0] _2078;
    wire [3:0] _2081;
    wire _2083;
    wire _2084;
    wire _3647;
    wire _3648;
    wire _3649;
    wire _3650;
    wire _150;
    reg _496;
    wire [3:0] _2040;
    wire [3:0] _2037;
    wire [3:0] _2034;
    wire [3:0] _2032;
    wire [3:0] _2035;
    wire [3:0] _2038;
    wire [3:0] _2041;
    wire [3:0] _2044;
    wire [3:0] _2047;
    wire [3:0] _2050;
    wire [3:0] _2053;
    wire _2055;
    wire _2056;
    wire _3651;
    wire _3652;
    wire _3653;
    wire _3654;
    wire _151;
    reg _501;
    wire [3:0] _2012;
    wire [3:0] _2009;
    wire [3:0] _2006;
    wire [3:0] _2004;
    wire [3:0] _2007;
    wire [3:0] _2010;
    wire [3:0] _2013;
    wire [3:0] _2016;
    wire [3:0] _2019;
    wire [3:0] _2022;
    wire [3:0] _2025;
    wire _2027;
    wire _2028;
    wire _3655;
    wire _3656;
    wire _3657;
    wire _3658;
    wire _152;
    reg _506;
    wire [3:0] _2255;
    wire [3:0] _2252;
    wire [3:0] _2249;
    wire [3:0] _2247;
    wire [3:0] _2250;
    wire [3:0] _2253;
    wire [3:0] _2256;
    wire [3:0] _2259;
    wire _2261;
    wire _2262;
    wire _3659;
    wire _3660;
    wire _3661;
    wire _3662;
    wire _153;
    reg _461;
    wire [3:0] _2520;
    wire [3:0] _2517;
    wire [3:0] _2514;
    wire [3:0] _2511;
    wire [3:0] _2509;
    wire [3:0] _2512;
    wire [3:0] _2515;
    wire [3:0] _2518;
    wire [3:0] _2521;
    wire _2523;
    wire _2524;
    wire _3663;
    wire _3664;
    wire _3665;
    wire _3666;
    wire _154;
    reg _411;
    wire [3:0] _2271;
    wire [3:0] _2268;
    wire [3:0] _2266;
    wire [3:0] _2269;
    wire [3:0] _2272;
    wire [3:0] _2275;
    wire [3:0] _2278;
    wire [3:0] _2281;
    wire [3:0] _2284;
    wire [3:0] _2287;
    wire _2289;
    wire _2290;
    wire _3667;
    wire _3668;
    wire _3669;
    wire _3670;
    wire _155;
    reg _456;
    wire [3:0] _2305;
    wire [3:0] _2302;
    wire [3:0] _2299;
    wire [3:0] _2296;
    wire [3:0] _2294;
    wire [3:0] _2297;
    wire [3:0] _2300;
    wire [3:0] _2303;
    wire [3:0] _2306;
    wire [3:0] _2309;
    wire [3:0] _2312;
    wire [3:0] _2315;
    wire _2317;
    wire _2318;
    wire _3671;
    wire _3672;
    wire _3673;
    wire _3674;
    wire _156;
    reg _451;
    wire [3:0] _2333;
    wire [3:0] _2330;
    wire [3:0] _2327;
    wire [3:0] _2324;
    wire [3:0] _2322;
    wire [3:0] _2325;
    wire [3:0] _2328;
    wire [3:0] _2331;
    wire [3:0] _2334;
    wire [3:0] _2337;
    wire [3:0] _2340;
    wire [3:0] _2343;
    wire _2345;
    wire _2346;
    wire _3675;
    wire _3676;
    wire _3677;
    wire _3678;
    wire _157;
    reg _446;
    wire [3:0] _2361;
    wire [3:0] _2358;
    wire [3:0] _2355;
    wire [3:0] _2352;
    wire [3:0] _2350;
    wire [3:0] _2353;
    wire [3:0] _2356;
    wire [3:0] _2359;
    wire [3:0] _2362;
    wire [3:0] _2365;
    wire [3:0] _2368;
    wire [3:0] _2371;
    wire _2373;
    wire _2374;
    wire _3679;
    wire _3680;
    wire _3681;
    wire _3682;
    wire _158;
    reg _441;
    wire [3:0] _2389;
    wire [3:0] _2386;
    wire [3:0] _2383;
    wire [3:0] _2380;
    wire [3:0] _2378;
    wire [3:0] _2381;
    wire [3:0] _2384;
    wire [3:0] _2387;
    wire [3:0] _2390;
    wire [3:0] _2393;
    wire [3:0] _2396;
    wire [3:0] _2399;
    wire _2401;
    wire _2402;
    wire _3683;
    wire _3684;
    wire _3685;
    wire _3686;
    wire _159;
    reg _436;
    wire [3:0] _2417;
    wire [3:0] _2414;
    wire [3:0] _2411;
    wire [3:0] _2408;
    wire [3:0] _2406;
    wire [3:0] _2409;
    wire [3:0] _2412;
    wire [3:0] _2415;
    wire [3:0] _2418;
    wire [3:0] _2421;
    wire [3:0] _2424;
    wire [3:0] _2427;
    wire _2429;
    wire _2430;
    wire _3687;
    wire _3688;
    wire _3689;
    wire _3690;
    wire _160;
    reg _431;
    wire [3:0] _2445;
    wire [3:0] _2442;
    wire [3:0] _2439;
    wire [3:0] _2436;
    wire [3:0] _2434;
    wire [3:0] _2437;
    wire [3:0] _2440;
    wire [3:0] _2443;
    wire [3:0] _2446;
    wire [3:0] _2449;
    wire [3:0] _2452;
    wire [3:0] _2455;
    wire _2457;
    wire _2458;
    wire _3691;
    wire _3692;
    wire _3693;
    wire _3694;
    wire _161;
    reg _426;
    wire [3:0] _2473;
    wire [3:0] _2470;
    wire [3:0] _2467;
    wire [3:0] _2464;
    wire [3:0] _2462;
    wire [3:0] _2465;
    wire [3:0] _2468;
    wire [3:0] _2471;
    wire [3:0] _2474;
    wire [3:0] _2477;
    wire [3:0] _2480;
    wire [3:0] _2483;
    wire _2485;
    wire _2486;
    wire _3695;
    wire _3696;
    wire _3697;
    wire _3698;
    wire _162;
    reg _421;
    wire [3:0] _2495;
    wire [3:0] _2492;
    wire [3:0] _2490;
    wire [3:0] _2493;
    wire [3:0] _2496;
    wire [3:0] _2499;
    wire [3:0] _2502;
    wire _2504;
    wire _2505;
    wire _3699;
    wire _3700;
    wire _3701;
    wire _3702;
    wire _163;
    reg _416;
    wire [3:0] _2760;
    wire [3:0] _2757;
    wire [3:0] _2754;
    wire [3:0] _2752;
    wire [3:0] _2755;
    wire [3:0] _2758;
    wire [3:0] _2761;
    wire [3:0] _2764;
    wire _2766;
    wire _2767;
    wire _3703;
    wire _3704;
    wire _3705;
    wire _3706;
    wire _164;
    reg _366;
    wire [3:0] _2732;
    wire [3:0] _2729;
    wire [3:0] _2726;
    wire [3:0] _2724;
    wire [3:0] _2727;
    wire [3:0] _2730;
    wire [3:0] _2733;
    wire [3:0] _2736;
    wire [3:0] _2739;
    wire [3:0] _2742;
    wire [3:0] _2745;
    wire _2747;
    wire _2748;
    wire _3707;
    wire _3708;
    wire _3709;
    wire _3710;
    wire _165;
    reg _371;
    wire [3:0] _2704;
    wire [3:0] _2701;
    wire [3:0] _2698;
    wire [3:0] _2696;
    wire [3:0] _2699;
    wire [3:0] _2702;
    wire [3:0] _2705;
    wire [3:0] _2708;
    wire [3:0] _2711;
    wire [3:0] _2714;
    wire [3:0] _2717;
    wire _2719;
    wire _2720;
    wire _3711;
    wire _3712;
    wire _3713;
    wire _3714;
    wire _166;
    reg _376;
    wire [3:0] _2676;
    wire [3:0] _2673;
    wire [3:0] _2670;
    wire [3:0] _2668;
    wire [3:0] _2671;
    wire [3:0] _2674;
    wire [3:0] _2677;
    wire [3:0] _2680;
    wire [3:0] _2683;
    wire [3:0] _2686;
    wire [3:0] _2689;
    wire _2691;
    wire _2692;
    wire _3715;
    wire _3716;
    wire _3717;
    wire _3718;
    wire _167;
    reg _381;
    wire [3:0] _2648;
    wire [3:0] _2645;
    wire [3:0] _2642;
    wire [3:0] _2640;
    wire [3:0] _2643;
    wire [3:0] _2646;
    wire [3:0] _2649;
    wire [3:0] _2652;
    wire [3:0] _2655;
    wire [3:0] _2658;
    wire [3:0] _2661;
    wire _2663;
    wire _2664;
    wire _3719;
    wire _3720;
    wire _3721;
    wire _3722;
    wire _168;
    reg _386;
    wire [3:0] _2620;
    wire [3:0] _2617;
    wire [3:0] _2614;
    wire [3:0] _2612;
    wire [3:0] _2615;
    wire [3:0] _2618;
    wire [3:0] _2621;
    wire [3:0] _2624;
    wire [3:0] _2627;
    wire [3:0] _2630;
    wire [3:0] _2633;
    wire _2635;
    wire _2636;
    wire _3723;
    wire _3724;
    wire _3725;
    wire _3726;
    wire _169;
    reg _391;
    wire [3:0] _2592;
    wire [3:0] _2589;
    wire [3:0] _2586;
    wire [3:0] _2584;
    wire [3:0] _2587;
    wire [3:0] _2590;
    wire [3:0] _2593;
    wire [3:0] _2596;
    wire [3:0] _2599;
    wire [3:0] _2602;
    wire [3:0] _2605;
    wire _2607;
    wire _2608;
    wire _3727;
    wire _3728;
    wire _3729;
    wire _3730;
    wire _170;
    reg _396;
    wire [3:0] _2564;
    wire [3:0] _2561;
    wire [3:0] _2558;
    wire [3:0] _2556;
    wire [3:0] _2559;
    wire [3:0] _2562;
    wire [3:0] _2565;
    wire [3:0] _2568;
    wire [3:0] _2571;
    wire [3:0] _2574;
    wire [3:0] _2577;
    wire _2579;
    wire _2580;
    wire _3731;
    wire _3732;
    wire _3733;
    wire _3734;
    wire _171;
    reg _401;
    wire [3:0] _2536;
    wire [3:0] _2533;
    wire [3:0] _2530;
    wire [3:0] _2528;
    wire [3:0] _2531;
    wire [3:0] _2534;
    wire [3:0] _2537;
    wire [3:0] _2540;
    wire [3:0] _2543;
    wire [3:0] _2546;
    wire [3:0] _2549;
    wire _2551;
    wire _2552;
    wire _3735;
    wire _3736;
    wire _3737;
    wire _3738;
    wire _172;
    reg _406;
    wire [3:0] _2779;
    wire [3:0] _2776;
    wire [3:0] _2773;
    wire [3:0] _2771;
    wire [3:0] _2774;
    wire [3:0] _2777;
    wire [3:0] _2780;
    wire [3:0] _2783;
    wire _2785;
    wire _2786;
    wire _3739;
    wire _3740;
    wire _3741;
    wire _3742;
    wire _173;
    reg _361;
    wire [3:0] _3044;
    wire [3:0] _3041;
    wire [3:0] _3038;
    wire [3:0] _3035;
    wire [3:0] _3033;
    wire [3:0] _3036;
    wire [3:0] _3039;
    wire [3:0] _3042;
    wire [3:0] _3045;
    wire _3047;
    wire _3048;
    wire _3743;
    wire _3744;
    wire _3745;
    wire _3746;
    wire _174;
    reg _311;
    wire [3:0] _2795;
    wire [3:0] _2792;
    wire [3:0] _2790;
    wire [3:0] _2793;
    wire [3:0] _2796;
    wire [3:0] _2799;
    wire [3:0] _2802;
    wire [3:0] _2805;
    wire [3:0] _2808;
    wire [3:0] _2811;
    wire _2813;
    wire _2814;
    wire _3747;
    wire _3748;
    wire _3749;
    wire _3750;
    wire _175;
    reg _356;
    wire [3:0] _2829;
    wire [3:0] _2826;
    wire [3:0] _2823;
    wire [3:0] _2820;
    wire [3:0] _2818;
    wire [3:0] _2821;
    wire [3:0] _2824;
    wire [3:0] _2827;
    wire [3:0] _2830;
    wire [3:0] _2833;
    wire [3:0] _2836;
    wire [3:0] _2839;
    wire _2841;
    wire _2842;
    wire _3751;
    wire _3752;
    wire _3753;
    wire _3754;
    wire _176;
    reg _351;
    wire [3:0] _2857;
    wire [3:0] _2854;
    wire [3:0] _2851;
    wire [3:0] _2848;
    wire [3:0] _2846;
    wire [3:0] _2849;
    wire [3:0] _2852;
    wire [3:0] _2855;
    wire [3:0] _2858;
    wire [3:0] _2861;
    wire [3:0] _2864;
    wire [3:0] _2867;
    wire _2869;
    wire _2870;
    wire _3755;
    wire _3756;
    wire _3757;
    wire _3758;
    wire _177;
    reg _346;
    wire [3:0] _2885;
    wire [3:0] _2882;
    wire [3:0] _2879;
    wire [3:0] _2876;
    wire [3:0] _2874;
    wire [3:0] _2877;
    wire [3:0] _2880;
    wire [3:0] _2883;
    wire [3:0] _2886;
    wire [3:0] _2889;
    wire [3:0] _2892;
    wire [3:0] _2895;
    wire _2897;
    wire _2898;
    wire _3759;
    wire _3760;
    wire _3761;
    wire _3762;
    wire _178;
    reg _341;
    wire [3:0] _2913;
    wire [3:0] _2910;
    wire [3:0] _2907;
    wire [3:0] _2904;
    wire [3:0] _2902;
    wire [3:0] _2905;
    wire [3:0] _2908;
    wire [3:0] _2911;
    wire [3:0] _2914;
    wire [3:0] _2917;
    wire [3:0] _2920;
    wire [3:0] _2923;
    wire _2925;
    wire _2926;
    wire _3763;
    wire _3764;
    wire _3765;
    wire _3766;
    wire _179;
    reg _336;
    wire [3:0] _2941;
    wire [3:0] _2938;
    wire [3:0] _2935;
    wire [3:0] _2932;
    wire [3:0] _2930;
    wire [3:0] _2933;
    wire [3:0] _2936;
    wire [3:0] _2939;
    wire [3:0] _2942;
    wire [3:0] _2945;
    wire [3:0] _2948;
    wire [3:0] _2951;
    wire _2953;
    wire _2954;
    wire _3767;
    wire _3768;
    wire _3769;
    wire _3770;
    wire _180;
    reg _331;
    wire [3:0] _2969;
    wire [3:0] _2966;
    wire [3:0] _2963;
    wire [3:0] _2960;
    wire [3:0] _2958;
    wire [3:0] _2961;
    wire [3:0] _2964;
    wire [3:0] _2967;
    wire [3:0] _2970;
    wire [3:0] _2973;
    wire [3:0] _2976;
    wire [3:0] _2979;
    wire _2981;
    wire _2982;
    wire _3771;
    wire _3772;
    wire _3773;
    wire _3774;
    wire _181;
    reg _326;
    wire [3:0] _2997;
    wire [3:0] _2994;
    wire [3:0] _2991;
    wire [3:0] _2988;
    wire [3:0] _2986;
    wire [3:0] _2989;
    wire [3:0] _2992;
    wire [3:0] _2995;
    wire [3:0] _2998;
    wire [3:0] _3001;
    wire [3:0] _3004;
    wire [3:0] _3007;
    wire _3009;
    wire _3010;
    wire _3775;
    wire _3776;
    wire _3777;
    wire _3778;
    wire _182;
    reg _321;
    wire [3:0] _3019;
    wire [3:0] _3016;
    wire [3:0] _3014;
    wire [3:0] _3017;
    wire [3:0] _3020;
    wire [3:0] _3023;
    wire [3:0] _3026;
    wire _3028;
    wire _3029;
    wire _3779;
    wire _3780;
    wire _3781;
    wire _3782;
    wire _183;
    reg _316;
    wire [3:0] _3284;
    wire [3:0] _3281;
    wire [3:0] _3278;
    wire [3:0] _3276;
    wire [3:0] _3279;
    wire [3:0] _3282;
    wire [3:0] _3285;
    wire [3:0] _3288;
    wire _3290;
    wire _3291;
    wire _3783;
    wire _3784;
    wire _3785;
    wire _3786;
    wire _184;
    reg _266;
    wire [3:0] _3256;
    wire [3:0] _3253;
    wire [3:0] _3250;
    wire [3:0] _3248;
    wire [3:0] _3251;
    wire [3:0] _3254;
    wire [3:0] _3257;
    wire [3:0] _3260;
    wire [3:0] _3263;
    wire [3:0] _3266;
    wire [3:0] _3269;
    wire _3271;
    wire _3272;
    wire _3787;
    wire _3788;
    wire _3789;
    wire _3790;
    wire _185;
    reg _271;
    wire [3:0] _3228;
    wire [3:0] _3225;
    wire [3:0] _3222;
    wire [3:0] _3220;
    wire [3:0] _3223;
    wire [3:0] _3226;
    wire [3:0] _3229;
    wire [3:0] _3232;
    wire [3:0] _3235;
    wire [3:0] _3238;
    wire [3:0] _3241;
    wire _3243;
    wire _3244;
    wire _3791;
    wire _3792;
    wire _3793;
    wire _3794;
    wire _186;
    reg _276;
    wire [3:0] _3200;
    wire [3:0] _3197;
    wire [3:0] _3194;
    wire [3:0] _3192;
    wire [3:0] _3195;
    wire [3:0] _3198;
    wire [3:0] _3201;
    wire [3:0] _3204;
    wire [3:0] _3207;
    wire [3:0] _3210;
    wire [3:0] _3213;
    wire _3215;
    wire _3216;
    wire _3795;
    wire _3796;
    wire _3797;
    wire _3798;
    wire _187;
    reg _281;
    wire [3:0] _3172;
    wire [3:0] _3169;
    wire [3:0] _3166;
    wire [3:0] _3164;
    wire [3:0] _3167;
    wire [3:0] _3170;
    wire [3:0] _3173;
    wire [3:0] _3176;
    wire [3:0] _3179;
    wire [3:0] _3182;
    wire [3:0] _3185;
    wire _3187;
    wire _3188;
    wire _3799;
    wire _3800;
    wire _3801;
    wire _3802;
    wire _188;
    reg _286;
    wire [3:0] _3144;
    wire [3:0] _3141;
    wire [3:0] _3138;
    wire [3:0] _3136;
    wire [3:0] _3139;
    wire [3:0] _3142;
    wire [3:0] _3145;
    wire [3:0] _3148;
    wire [3:0] _3151;
    wire [3:0] _3154;
    wire [3:0] _3157;
    wire _3159;
    wire _3160;
    wire _3803;
    wire _3804;
    wire _3805;
    wire _3806;
    wire _189;
    reg _291;
    wire [3:0] _3116;
    wire [3:0] _3113;
    wire [3:0] _3110;
    wire [3:0] _3108;
    wire [3:0] _3111;
    wire [3:0] _3114;
    wire [3:0] _3117;
    wire [3:0] _3120;
    wire [3:0] _3123;
    wire [3:0] _3126;
    wire [3:0] _3129;
    wire _3131;
    wire _3132;
    wire _3807;
    wire _3808;
    wire _3809;
    wire _3810;
    wire _190;
    reg _296;
    wire [3:0] _3088;
    wire [3:0] _3085;
    wire [3:0] _3082;
    wire [3:0] _3080;
    wire [3:0] _3083;
    wire [3:0] _3086;
    wire [3:0] _3089;
    wire [3:0] _3092;
    wire [3:0] _3095;
    wire [3:0] _3098;
    wire [3:0] _3101;
    wire _3103;
    wire _3104;
    wire _3811;
    wire _3812;
    wire _3813;
    wire _3814;
    wire _191;
    reg _301;
    wire [3:0] _3060;
    wire [3:0] _3057;
    wire [3:0] _3054;
    wire [3:0] _3052;
    wire [3:0] _3055;
    wire [3:0] _3058;
    wire [3:0] _3061;
    wire [3:0] _3064;
    wire [3:0] _3067;
    wire [3:0] _3070;
    wire [3:0] _3073;
    wire _3075;
    wire _3076;
    wire _3815;
    wire _3816;
    wire _3817;
    wire _3818;
    wire _192;
    reg _306;
    wire [3:0] _3297;
    wire [3:0] _3295;
    wire [3:0] _3298;
    wire [3:0] _3301;
    wire _3303;
    wire _3304;
    wire _3819;
    wire _3820;
    wire _3821;
    wire _3822;
    wire _193;
    reg _261;
    wire [3:0] _3310;
    wire [3:0] _3308;
    wire [3:0] _3311;
    wire [3:0] _3314;
    wire [3:0] _3317;
    wire [3:0] _3320;
    wire _3322;
    wire _3323;
    wire _3823;
    wire _3824;
    wire _3825;
    wire _3826;
    wire _194;
    reg _256;
    wire [3:0] _3329;
    wire [3:0] _3327;
    wire [3:0] _3330;
    wire [3:0] _3333;
    wire [3:0] _3336;
    wire [3:0] _3339;
    wire _3341;
    wire _3342;
    wire _3827;
    wire _3828;
    wire _3829;
    wire _3830;
    wire _195;
    reg _251;
    wire [3:0] _3348;
    wire [3:0] _3346;
    wire [3:0] _3349;
    wire [3:0] _3352;
    wire [3:0] _3355;
    wire [3:0] _3358;
    wire _3360;
    wire _3361;
    wire _3831;
    wire _3832;
    wire _3833;
    wire _3834;
    wire _196;
    reg _246;
    wire [3:0] _3367;
    wire [3:0] _3365;
    wire [3:0] _3368;
    wire [3:0] _3371;
    wire [3:0] _3374;
    wire [3:0] _3377;
    wire _3379;
    wire _3380;
    wire _3835;
    wire _3836;
    wire _3837;
    wire _3838;
    wire _197;
    reg _241;
    wire [3:0] _3386;
    wire [3:0] _3384;
    wire [3:0] _3387;
    wire [3:0] _3390;
    wire [3:0] _3393;
    wire [3:0] _3396;
    wire _3398;
    wire _3399;
    wire _3839;
    wire _3840;
    wire _3841;
    wire _3842;
    wire _198;
    reg _236;
    wire [3:0] _3405;
    wire [3:0] _3403;
    wire [3:0] _3406;
    wire [3:0] _3409;
    wire [3:0] _3412;
    wire [3:0] _3415;
    wire _3417;
    wire _3418;
    wire _3843;
    wire _3844;
    wire _3845;
    wire _3846;
    wire _199;
    reg _231;
    wire [3:0] _3424;
    wire [3:0] _3422;
    wire [3:0] _3425;
    wire [3:0] _3428;
    wire [3:0] _3431;
    wire [3:0] _3434;
    wire _3436;
    wire _3437;
    wire _3847;
    wire _3848;
    wire _3849;
    wire _3850;
    wire _200;
    reg _226;
    wire [3:0] _3443;
    wire [3:0] _3441;
    wire [3:0] _3444;
    wire [3:0] _3447;
    wire [3:0] _3450;
    wire [3:0] _3453;
    wire _3455;
    wire _3456;
    wire _3851;
    wire _3852;
    wire _3853;
    wire _3854;
    wire _201;
    reg _221;
    wire [3:0] _3856;
    wire [3:0] _3859;
    wire [3:0] _3862;
    wire _3864;
    wire _203;
    wire _205;
    wire _207;
    wire _3866;
    wire _3867;
    wire _3868;
    wire _3869;
    wire _208;
    reg _217;
    wire _3865;
    wire gnd;
    wire _3870;
    wire _210;
    wire _3871;
    wire _211;
    wire [15:0] _719;
    wire [15:0] _722;
    wire [15:0] _725;
    wire [15:0] _728;
    wire [15:0] _731;
    wire [15:0] _734;
    wire [15:0] _737;
    wire [15:0] _740;
    wire [15:0] _743;
    wire [15:0] _746;
    wire [15:0] _749;
    wire [15:0] _752;
    wire [15:0] _755;
    wire [15:0] _758;
    wire [15:0] _761;
    wire [15:0] _764;
    wire [15:0] _767;
    wire [15:0] _770;
    wire [15:0] _773;
    wire [15:0] _776;
    wire [15:0] _779;
    wire [15:0] _782;
    wire [15:0] _785;
    wire [15:0] _788;
    wire [15:0] _791;
    wire [15:0] _794;
    wire [15:0] _797;
    wire [15:0] _800;
    wire [15:0] _803;
    wire [15:0] _806;
    wire [15:0] _809;
    wire [15:0] _812;
    wire [15:0] _815;
    wire [15:0] _818;
    wire [15:0] _821;
    wire [15:0] _824;
    wire [15:0] _827;
    wire [15:0] _830;
    wire [15:0] _833;
    wire [15:0] _836;
    wire [15:0] _839;
    wire [15:0] _842;
    wire [15:0] _845;
    wire [15:0] _848;
    wire [15:0] _851;
    wire [15:0] _854;
    wire [15:0] _857;
    wire [15:0] _860;
    wire [15:0] _863;
    wire [15:0] _866;
    wire [15:0] _869;
    wire [15:0] _872;
    wire [15:0] _875;
    wire [15:0] _878;
    wire [15:0] _881;
    wire [15:0] _884;
    wire [15:0] _887;
    wire [15:0] _890;
    wire [15:0] _893;
    wire [15:0] _896;
    wire [15:0] _899;
    wire [15:0] _902;
    wire [15:0] _905;
    wire [15:0] _908;
    wire [15:0] _911;
    wire [15:0] _914;
    wire [15:0] _917;
    wire [15:0] _920;
    wire [15:0] _923;
    wire [15:0] _926;
    wire [15:0] _929;
    wire [15:0] _932;
    wire [15:0] _935;
    wire [15:0] _938;
    wire [15:0] _941;
    wire [15:0] _944;
    wire [15:0] _947;
    wire [15:0] _950;
    wire [15:0] _953;
    wire [15:0] _956;
    wire [15:0] _959;
    wire [15:0] _962;
    wire [15:0] _965;
    wire [15:0] _968;
    wire [15:0] _971;
    wire [15:0] _974;
    wire [15:0] _977;
    wire [15:0] _980;
    wire [15:0] _983;
    wire [15:0] _986;
    wire [15:0] _989;
    wire [15:0] _992;
    wire [15:0] _995;
    wire [15:0] _998;
    wire [15:0] _1001;
    wire [15:0] _1004;
    wire [15:0] _1007;
    wire [15:0] _1010;
    wire [15:0] _1013;
    wire [15:0] _1016;
    wire _3873;
    wire _213;
    wire _3874;
    assign _709 = 15'b000000000000000;
    assign _712 = { _709,
                    _711 };
    assign _707 = { _709,
                    _706 };
    assign _702 = { _709,
                    _701 };
    assign _697 = { _709,
                    _696 };
    assign _692 = { _709,
                    _691 };
    assign _687 = { _709,
                    _686 };
    assign _682 = { _709,
                    _681 };
    assign _677 = { _709,
                    _676 };
    assign _672 = { _709,
                    _671 };
    assign _667 = { _709,
                    _666 };
    assign _662 = { _709,
                    _661 };
    assign _657 = { _709,
                    _656 };
    assign _652 = { _709,
                    _651 };
    assign _647 = { _709,
                    _646 };
    assign _642 = { _709,
                    _641 };
    assign _637 = { _709,
                    _636 };
    assign _632 = { _709,
                    _631 };
    assign _627 = { _709,
                    _626 };
    assign _622 = { _709,
                    _621 };
    assign _617 = { _709,
                    _616 };
    assign _612 = { _709,
                    _611 };
    assign _607 = { _709,
                    _606 };
    assign _602 = { _709,
                    _601 };
    assign _597 = { _709,
                    _596 };
    assign _592 = { _709,
                    _591 };
    assign _587 = { _709,
                    _586 };
    assign _582 = { _709,
                    _581 };
    assign _577 = { _709,
                    _576 };
    assign _572 = { _709,
                    _571 };
    assign _567 = { _709,
                    _566 };
    assign _562 = { _709,
                    _561 };
    assign _557 = { _709,
                    _556 };
    assign _552 = { _709,
                    _551 };
    assign _547 = { _709,
                    _546 };
    assign _542 = { _709,
                    _541 };
    assign _537 = { _709,
                    _536 };
    assign _532 = { _709,
                    _531 };
    assign _527 = { _709,
                    _526 };
    assign _522 = { _709,
                    _521 };
    assign _517 = { _709,
                    _516 };
    assign _512 = { _709,
                    _511 };
    assign _507 = { _709,
                    _506 };
    assign _502 = { _709,
                    _501 };
    assign _497 = { _709,
                    _496 };
    assign _492 = { _709,
                    _491 };
    assign _487 = { _709,
                    _486 };
    assign _482 = { _709,
                    _481 };
    assign _477 = { _709,
                    _476 };
    assign _472 = { _709,
                    _471 };
    assign _467 = { _709,
                    _466 };
    assign _462 = { _709,
                    _461 };
    assign _457 = { _709,
                    _456 };
    assign _452 = { _709,
                    _451 };
    assign _447 = { _709,
                    _446 };
    assign _442 = { _709,
                    _441 };
    assign _437 = { _709,
                    _436 };
    assign _432 = { _709,
                    _431 };
    assign _427 = { _709,
                    _426 };
    assign _422 = { _709,
                    _421 };
    assign _417 = { _709,
                    _416 };
    assign _412 = { _709,
                    _411 };
    assign _407 = { _709,
                    _406 };
    assign _402 = { _709,
                    _401 };
    assign _397 = { _709,
                    _396 };
    assign _392 = { _709,
                    _391 };
    assign _387 = { _709,
                    _386 };
    assign _382 = { _709,
                    _381 };
    assign _377 = { _709,
                    _376 };
    assign _372 = { _709,
                    _371 };
    assign _367 = { _709,
                    _366 };
    assign _362 = { _709,
                    _361 };
    assign _357 = { _709,
                    _356 };
    assign _352 = { _709,
                    _351 };
    assign _347 = { _709,
                    _346 };
    assign _342 = { _709,
                    _341 };
    assign _337 = { _709,
                    _336 };
    assign _332 = { _709,
                    _331 };
    assign _327 = { _709,
                    _326 };
    assign _322 = { _709,
                    _321 };
    assign _317 = { _709,
                    _316 };
    assign _312 = { _709,
                    _311 };
    assign _307 = { _709,
                    _306 };
    assign _302 = { _709,
                    _301 };
    assign _297 = { _709,
                    _296 };
    assign _292 = { _709,
                    _291 };
    assign _287 = { _709,
                    _286 };
    assign _282 = { _709,
                    _281 };
    assign _277 = { _709,
                    _276 };
    assign _272 = { _709,
                    _271 };
    assign _267 = { _709,
                    _266 };
    assign _262 = { _709,
                    _261 };
    assign _257 = { _709,
                    _256 };
    assign _252 = { _709,
                    _251 };
    assign _247 = { _709,
                    _246 };
    assign _242 = { _709,
                    _241 };
    assign _237 = { _709,
                    _236 };
    assign _232 = { _709,
                    _231 };
    assign _227 = { _709,
                    _226 };
    assign _222 = { _709,
                    _221 };
    assign _218 = { _709,
                    _217 };
    assign _223 = _218 + _222;
    assign _228 = _223 + _227;
    assign _233 = _228 + _232;
    assign _238 = _233 + _237;
    assign _243 = _238 + _242;
    assign _248 = _243 + _247;
    assign _253 = _248 + _252;
    assign _258 = _253 + _257;
    assign _263 = _258 + _262;
    assign _268 = _263 + _267;
    assign _273 = _268 + _272;
    assign _278 = _273 + _277;
    assign _283 = _278 + _282;
    assign _288 = _283 + _287;
    assign _293 = _288 + _292;
    assign _298 = _293 + _297;
    assign _303 = _298 + _302;
    assign _308 = _303 + _307;
    assign _313 = _308 + _312;
    assign _318 = _313 + _317;
    assign _323 = _318 + _322;
    assign _328 = _323 + _327;
    assign _333 = _328 + _332;
    assign _338 = _333 + _337;
    assign _343 = _338 + _342;
    assign _348 = _343 + _347;
    assign _353 = _348 + _352;
    assign _358 = _353 + _357;
    assign _363 = _358 + _362;
    assign _368 = _363 + _367;
    assign _373 = _368 + _372;
    assign _378 = _373 + _377;
    assign _383 = _378 + _382;
    assign _388 = _383 + _387;
    assign _393 = _388 + _392;
    assign _398 = _393 + _397;
    assign _403 = _398 + _402;
    assign _408 = _403 + _407;
    assign _413 = _408 + _412;
    assign _418 = _413 + _417;
    assign _423 = _418 + _422;
    assign _428 = _423 + _427;
    assign _433 = _428 + _432;
    assign _438 = _433 + _437;
    assign _443 = _438 + _442;
    assign _448 = _443 + _447;
    assign _453 = _448 + _452;
    assign _458 = _453 + _457;
    assign _463 = _458 + _462;
    assign _468 = _463 + _467;
    assign _473 = _468 + _472;
    assign _478 = _473 + _477;
    assign _483 = _478 + _482;
    assign _488 = _483 + _487;
    assign _493 = _488 + _492;
    assign _498 = _493 + _497;
    assign _503 = _498 + _502;
    assign _508 = _503 + _507;
    assign _513 = _508 + _512;
    assign _518 = _513 + _517;
    assign _523 = _518 + _522;
    assign _528 = _523 + _527;
    assign _533 = _528 + _532;
    assign _538 = _533 + _537;
    assign _543 = _538 + _542;
    assign _548 = _543 + _547;
    assign _553 = _548 + _552;
    assign _558 = _553 + _557;
    assign _563 = _558 + _562;
    assign _568 = _563 + _567;
    assign _573 = _568 + _572;
    assign _578 = _573 + _577;
    assign _583 = _578 + _582;
    assign _588 = _583 + _587;
    assign _593 = _588 + _592;
    assign _598 = _593 + _597;
    assign _603 = _598 + _602;
    assign _608 = _603 + _607;
    assign _613 = _608 + _612;
    assign _618 = _613 + _617;
    assign _623 = _618 + _622;
    assign _628 = _623 + _627;
    assign _633 = _628 + _632;
    assign _638 = _633 + _637;
    assign _643 = _638 + _642;
    assign _648 = _643 + _647;
    assign _653 = _648 + _652;
    assign _658 = _653 + _657;
    assign _663 = _658 + _662;
    assign _668 = _663 + _667;
    assign _673 = _668 + _672;
    assign _678 = _673 + _677;
    assign _683 = _678 + _682;
    assign _688 = _683 + _687;
    assign _693 = _688 + _692;
    assign _698 = _693 + _697;
    assign _703 = _698 + _702;
    assign _708 = _703 + _707;
    assign _713 = _708 + _712;
    assign _714 = 16'b0000000000000000;
    assign _1017 = _715 + _1016;
    assign _717 = _203 ? _714 : _715;
    assign _1018 = _213 ? _1017 : _717;
    assign _2 = _1018;
    always @(posedge _205) begin
        if (_203)
            _715 <= _714;
        else
            _715 <= _2;
    end
    assign _1031 = _213 ? _1030 : gnd;
    assign _1032 = _210 ? gnd : _1031;
    assign _4 = _1032;
    assign _1015 = { _709,
                     _4 };
    assign _1050 = _213 ? _1049 : gnd;
    assign _1051 = _210 ? gnd : _1050;
    assign _5 = _1051;
    assign _1012 = { _709,
                     _5 };
    assign _1069 = _213 ? _1068 : gnd;
    assign _1070 = _210 ? gnd : _1069;
    assign _6 = _1070;
    assign _1009 = { _709,
                     _6 };
    assign _1088 = _213 ? _1087 : gnd;
    assign _1089 = _210 ? gnd : _1088;
    assign _7 = _1089;
    assign _1006 = { _709,
                     _7 };
    assign _1107 = _213 ? _1106 : gnd;
    assign _1108 = _210 ? gnd : _1107;
    assign _8 = _1108;
    assign _1003 = { _709,
                     _8 };
    assign _1126 = _213 ? _1125 : gnd;
    assign _1127 = _210 ? gnd : _1126;
    assign _9 = _1127;
    assign _1000 = { _709,
                     _9 };
    assign _1145 = _213 ? _1144 : gnd;
    assign _1146 = _210 ? gnd : _1145;
    assign _10 = _1146;
    assign _997 = { _709,
                    _10 };
    assign _1164 = _213 ? _1163 : gnd;
    assign _1165 = _210 ? gnd : _1164;
    assign _11 = _1165;
    assign _994 = { _709,
                    _11 };
    assign _1183 = _213 ? _1182 : gnd;
    assign _1184 = _210 ? gnd : _1183;
    assign _12 = _1184;
    assign _991 = { _709,
                    _12 };
    assign _1196 = _213 ? _1195 : gnd;
    assign _1197 = _210 ? gnd : _1196;
    assign _13 = _1197;
    assign _988 = { _709,
                    _13 };
    assign _1215 = _213 ? _1214 : gnd;
    assign _1216 = _210 ? gnd : _1215;
    assign _14 = _1216;
    assign _985 = { _709,
                    _14 };
    assign _1243 = _213 ? _1242 : gnd;
    assign _1244 = _210 ? gnd : _1243;
    assign _15 = _1244;
    assign _982 = { _709,
                    _15 };
    assign _1271 = _213 ? _1270 : gnd;
    assign _1272 = _210 ? gnd : _1271;
    assign _16 = _1272;
    assign _979 = { _709,
                    _16 };
    assign _1299 = _213 ? _1298 : gnd;
    assign _1300 = _210 ? gnd : _1299;
    assign _17 = _1300;
    assign _976 = { _709,
                    _17 };
    assign _1327 = _213 ? _1326 : gnd;
    assign _1328 = _210 ? gnd : _1327;
    assign _18 = _1328;
    assign _973 = { _709,
                    _18 };
    assign _1355 = _213 ? _1354 : gnd;
    assign _1356 = _210 ? gnd : _1355;
    assign _19 = _1356;
    assign _970 = { _709,
                    _19 };
    assign _1383 = _213 ? _1382 : gnd;
    assign _1384 = _210 ? gnd : _1383;
    assign _20 = _1384;
    assign _967 = { _709,
                    _20 };
    assign _1411 = _213 ? _1410 : gnd;
    assign _1412 = _210 ? gnd : _1411;
    assign _21 = _1412;
    assign _964 = { _709,
                    _21 };
    assign _1439 = _213 ? _1438 : gnd;
    assign _1440 = _210 ? gnd : _1439;
    assign _22 = _1440;
    assign _961 = { _709,
                    _22 };
    assign _1458 = _213 ? _1457 : gnd;
    assign _1459 = _210 ? gnd : _1458;
    assign _23 = _1459;
    assign _958 = { _709,
                    _23 };
    assign _1477 = _213 ? _1476 : gnd;
    assign _1478 = _210 ? gnd : _1477;
    assign _24 = _1478;
    assign _955 = { _709,
                    _24 };
    assign _1505 = _213 ? _1504 : gnd;
    assign _1506 = _210 ? gnd : _1505;
    assign _25 = _1506;
    assign _952 = { _709,
                    _25 };
    assign _1533 = _213 ? _1532 : gnd;
    assign _1534 = _210 ? gnd : _1533;
    assign _26 = _1534;
    assign _949 = { _709,
                    _26 };
    assign _1561 = _213 ? _1560 : gnd;
    assign _1562 = _210 ? gnd : _1561;
    assign _27 = _1562;
    assign _946 = { _709,
                    _27 };
    assign _1589 = _213 ? _1588 : gnd;
    assign _1590 = _210 ? gnd : _1589;
    assign _28 = _1590;
    assign _943 = { _709,
                    _28 };
    assign _1617 = _213 ? _1616 : gnd;
    assign _1618 = _210 ? gnd : _1617;
    assign _29 = _1618;
    assign _940 = { _709,
                    _29 };
    assign _1645 = _213 ? _1644 : gnd;
    assign _1646 = _210 ? gnd : _1645;
    assign _30 = _1646;
    assign _937 = { _709,
                    _30 };
    assign _1673 = _213 ? _1672 : gnd;
    assign _1674 = _210 ? gnd : _1673;
    assign _31 = _1674;
    assign _934 = { _709,
                    _31 };
    assign _1701 = _213 ? _1700 : gnd;
    assign _1702 = _210 ? gnd : _1701;
    assign _32 = _1702;
    assign _931 = { _709,
                    _32 };
    assign _1720 = _213 ? _1719 : gnd;
    assign _1721 = _210 ? gnd : _1720;
    assign _33 = _1721;
    assign _928 = { _709,
                    _33 };
    assign _1739 = _213 ? _1738 : gnd;
    assign _1740 = _210 ? gnd : _1739;
    assign _34 = _1740;
    assign _925 = { _709,
                    _34 };
    assign _1767 = _213 ? _1766 : gnd;
    assign _1768 = _210 ? gnd : _1767;
    assign _35 = _1768;
    assign _922 = { _709,
                    _35 };
    assign _1795 = _213 ? _1794 : gnd;
    assign _1796 = _210 ? gnd : _1795;
    assign _36 = _1796;
    assign _919 = { _709,
                    _36 };
    assign _1823 = _213 ? _1822 : gnd;
    assign _1824 = _210 ? gnd : _1823;
    assign _37 = _1824;
    assign _916 = { _709,
                    _37 };
    assign _1851 = _213 ? _1850 : gnd;
    assign _1852 = _210 ? gnd : _1851;
    assign _38 = _1852;
    assign _913 = { _709,
                    _38 };
    assign _1879 = _213 ? _1878 : gnd;
    assign _1880 = _210 ? gnd : _1879;
    assign _39 = _1880;
    assign _910 = { _709,
                    _39 };
    assign _1907 = _213 ? _1906 : gnd;
    assign _1908 = _210 ? gnd : _1907;
    assign _40 = _1908;
    assign _907 = { _709,
                    _40 };
    assign _1935 = _213 ? _1934 : gnd;
    assign _1936 = _210 ? gnd : _1935;
    assign _41 = _1936;
    assign _904 = { _709,
                    _41 };
    assign _1963 = _213 ? _1962 : gnd;
    assign _1964 = _210 ? gnd : _1963;
    assign _42 = _1964;
    assign _901 = { _709,
                    _42 };
    assign _1982 = _213 ? _1981 : gnd;
    assign _1983 = _210 ? gnd : _1982;
    assign _43 = _1983;
    assign _898 = { _709,
                    _43 };
    assign _2001 = _213 ? _2000 : gnd;
    assign _2002 = _210 ? gnd : _2001;
    assign _44 = _2002;
    assign _895 = { _709,
                    _44 };
    assign _2029 = _213 ? _2028 : gnd;
    assign _2030 = _210 ? gnd : _2029;
    assign _45 = _2030;
    assign _892 = { _709,
                    _45 };
    assign _2057 = _213 ? _2056 : gnd;
    assign _2058 = _210 ? gnd : _2057;
    assign _46 = _2058;
    assign _889 = { _709,
                    _46 };
    assign _2085 = _213 ? _2084 : gnd;
    assign _2086 = _210 ? gnd : _2085;
    assign _47 = _2086;
    assign _886 = { _709,
                    _47 };
    assign _2113 = _213 ? _2112 : gnd;
    assign _2114 = _210 ? gnd : _2113;
    assign _48 = _2114;
    assign _883 = { _709,
                    _48 };
    assign _2141 = _213 ? _2140 : gnd;
    assign _2142 = _210 ? gnd : _2141;
    assign _49 = _2142;
    assign _880 = { _709,
                    _49 };
    assign _2169 = _213 ? _2168 : gnd;
    assign _2170 = _210 ? gnd : _2169;
    assign _50 = _2170;
    assign _877 = { _709,
                    _50 };
    assign _2197 = _213 ? _2196 : gnd;
    assign _2198 = _210 ? gnd : _2197;
    assign _51 = _2198;
    assign _874 = { _709,
                    _51 };
    assign _2225 = _213 ? _2224 : gnd;
    assign _2226 = _210 ? gnd : _2225;
    assign _52 = _2226;
    assign _871 = { _709,
                    _52 };
    assign _2244 = _213 ? _2243 : gnd;
    assign _2245 = _210 ? gnd : _2244;
    assign _53 = _2245;
    assign _868 = { _709,
                    _53 };
    assign _2263 = _213 ? _2262 : gnd;
    assign _2264 = _210 ? gnd : _2263;
    assign _54 = _2264;
    assign _865 = { _709,
                    _54 };
    assign _2291 = _213 ? _2290 : gnd;
    assign _2292 = _210 ? gnd : _2291;
    assign _55 = _2292;
    assign _862 = { _709,
                    _55 };
    assign _2319 = _213 ? _2318 : gnd;
    assign _2320 = _210 ? gnd : _2319;
    assign _56 = _2320;
    assign _859 = { _709,
                    _56 };
    assign _2347 = _213 ? _2346 : gnd;
    assign _2348 = _210 ? gnd : _2347;
    assign _57 = _2348;
    assign _856 = { _709,
                    _57 };
    assign _2375 = _213 ? _2374 : gnd;
    assign _2376 = _210 ? gnd : _2375;
    assign _58 = _2376;
    assign _853 = { _709,
                    _58 };
    assign _2403 = _213 ? _2402 : gnd;
    assign _2404 = _210 ? gnd : _2403;
    assign _59 = _2404;
    assign _850 = { _709,
                    _59 };
    assign _2431 = _213 ? _2430 : gnd;
    assign _2432 = _210 ? gnd : _2431;
    assign _60 = _2432;
    assign _847 = { _709,
                    _60 };
    assign _2459 = _213 ? _2458 : gnd;
    assign _2460 = _210 ? gnd : _2459;
    assign _61 = _2460;
    assign _844 = { _709,
                    _61 };
    assign _2487 = _213 ? _2486 : gnd;
    assign _2488 = _210 ? gnd : _2487;
    assign _62 = _2488;
    assign _841 = { _709,
                    _62 };
    assign _2506 = _213 ? _2505 : gnd;
    assign _2507 = _210 ? gnd : _2506;
    assign _63 = _2507;
    assign _838 = { _709,
                    _63 };
    assign _2525 = _213 ? _2524 : gnd;
    assign _2526 = _210 ? gnd : _2525;
    assign _64 = _2526;
    assign _835 = { _709,
                    _64 };
    assign _2553 = _213 ? _2552 : gnd;
    assign _2554 = _210 ? gnd : _2553;
    assign _65 = _2554;
    assign _832 = { _709,
                    _65 };
    assign _2581 = _213 ? _2580 : gnd;
    assign _2582 = _210 ? gnd : _2581;
    assign _66 = _2582;
    assign _829 = { _709,
                    _66 };
    assign _2609 = _213 ? _2608 : gnd;
    assign _2610 = _210 ? gnd : _2609;
    assign _67 = _2610;
    assign _826 = { _709,
                    _67 };
    assign _2637 = _213 ? _2636 : gnd;
    assign _2638 = _210 ? gnd : _2637;
    assign _68 = _2638;
    assign _823 = { _709,
                    _68 };
    assign _2665 = _213 ? _2664 : gnd;
    assign _2666 = _210 ? gnd : _2665;
    assign _69 = _2666;
    assign _820 = { _709,
                    _69 };
    assign _2693 = _213 ? _2692 : gnd;
    assign _2694 = _210 ? gnd : _2693;
    assign _70 = _2694;
    assign _817 = { _709,
                    _70 };
    assign _2721 = _213 ? _2720 : gnd;
    assign _2722 = _210 ? gnd : _2721;
    assign _71 = _2722;
    assign _814 = { _709,
                    _71 };
    assign _2749 = _213 ? _2748 : gnd;
    assign _2750 = _210 ? gnd : _2749;
    assign _72 = _2750;
    assign _811 = { _709,
                    _72 };
    assign _2768 = _213 ? _2767 : gnd;
    assign _2769 = _210 ? gnd : _2768;
    assign _73 = _2769;
    assign _808 = { _709,
                    _73 };
    assign _2787 = _213 ? _2786 : gnd;
    assign _2788 = _210 ? gnd : _2787;
    assign _74 = _2788;
    assign _805 = { _709,
                    _74 };
    assign _2815 = _213 ? _2814 : gnd;
    assign _2816 = _210 ? gnd : _2815;
    assign _75 = _2816;
    assign _802 = { _709,
                    _75 };
    assign _2843 = _213 ? _2842 : gnd;
    assign _2844 = _210 ? gnd : _2843;
    assign _76 = _2844;
    assign _799 = { _709,
                    _76 };
    assign _2871 = _213 ? _2870 : gnd;
    assign _2872 = _210 ? gnd : _2871;
    assign _77 = _2872;
    assign _796 = { _709,
                    _77 };
    assign _2899 = _213 ? _2898 : gnd;
    assign _2900 = _210 ? gnd : _2899;
    assign _78 = _2900;
    assign _793 = { _709,
                    _78 };
    assign _2927 = _213 ? _2926 : gnd;
    assign _2928 = _210 ? gnd : _2927;
    assign _79 = _2928;
    assign _790 = { _709,
                    _79 };
    assign _2955 = _213 ? _2954 : gnd;
    assign _2956 = _210 ? gnd : _2955;
    assign _80 = _2956;
    assign _787 = { _709,
                    _80 };
    assign _2983 = _213 ? _2982 : gnd;
    assign _2984 = _210 ? gnd : _2983;
    assign _81 = _2984;
    assign _784 = { _709,
                    _81 };
    assign _3011 = _213 ? _3010 : gnd;
    assign _3012 = _210 ? gnd : _3011;
    assign _82 = _3012;
    assign _781 = { _709,
                    _82 };
    assign _3030 = _213 ? _3029 : gnd;
    assign _3031 = _210 ? gnd : _3030;
    assign _83 = _3031;
    assign _778 = { _709,
                    _83 };
    assign _3049 = _213 ? _3048 : gnd;
    assign _3050 = _210 ? gnd : _3049;
    assign _84 = _3050;
    assign _775 = { _709,
                    _84 };
    assign _3077 = _213 ? _3076 : gnd;
    assign _3078 = _210 ? gnd : _3077;
    assign _85 = _3078;
    assign _772 = { _709,
                    _85 };
    assign _3105 = _213 ? _3104 : gnd;
    assign _3106 = _210 ? gnd : _3105;
    assign _86 = _3106;
    assign _769 = { _709,
                    _86 };
    assign _3133 = _213 ? _3132 : gnd;
    assign _3134 = _210 ? gnd : _3133;
    assign _87 = _3134;
    assign _766 = { _709,
                    _87 };
    assign _3161 = _213 ? _3160 : gnd;
    assign _3162 = _210 ? gnd : _3161;
    assign _88 = _3162;
    assign _763 = { _709,
                    _88 };
    assign _3189 = _213 ? _3188 : gnd;
    assign _3190 = _210 ? gnd : _3189;
    assign _89 = _3190;
    assign _760 = { _709,
                    _89 };
    assign _3217 = _213 ? _3216 : gnd;
    assign _3218 = _210 ? gnd : _3217;
    assign _90 = _3218;
    assign _757 = { _709,
                    _90 };
    assign _3245 = _213 ? _3244 : gnd;
    assign _3246 = _210 ? gnd : _3245;
    assign _91 = _3246;
    assign _754 = { _709,
                    _91 };
    assign _3273 = _213 ? _3272 : gnd;
    assign _3274 = _210 ? gnd : _3273;
    assign _92 = _3274;
    assign _751 = { _709,
                    _92 };
    assign _3292 = _213 ? _3291 : gnd;
    assign _3293 = _210 ? gnd : _3292;
    assign _93 = _3293;
    assign _748 = { _709,
                    _93 };
    assign _3305 = _213 ? _3304 : gnd;
    assign _3306 = _210 ? gnd : _3305;
    assign _94 = _3306;
    assign _745 = { _709,
                    _94 };
    assign _3324 = _213 ? _3323 : gnd;
    assign _3325 = _210 ? gnd : _3324;
    assign _95 = _3325;
    assign _742 = { _709,
                    _95 };
    assign _3343 = _213 ? _3342 : gnd;
    assign _3344 = _210 ? gnd : _3343;
    assign _96 = _3344;
    assign _739 = { _709,
                    _96 };
    assign _3362 = _213 ? _3361 : gnd;
    assign _3363 = _210 ? gnd : _3362;
    assign _97 = _3363;
    assign _736 = { _709,
                    _97 };
    assign _3381 = _213 ? _3380 : gnd;
    assign _3382 = _210 ? gnd : _3381;
    assign _98 = _3382;
    assign _733 = { _709,
                    _98 };
    assign _3400 = _213 ? _3399 : gnd;
    assign _3401 = _210 ? gnd : _3400;
    assign _99 = _3401;
    assign _730 = { _709,
                    _99 };
    assign _3419 = _213 ? _3418 : gnd;
    assign _3420 = _210 ? gnd : _3419;
    assign _100 = _3420;
    assign _727 = { _709,
                    _100 };
    assign _3438 = _213 ? _3437 : gnd;
    assign _3439 = _210 ? gnd : _3438;
    assign _101 = _3439;
    assign _724 = { _709,
                    _101 };
    assign _3457 = _213 ? _3456 : gnd;
    assign _3458 = _210 ? gnd : _3457;
    assign _102 = _3458;
    assign _721 = { _709,
                    _102 };
    assign _3863 = 4'b0100;
    assign _3860 = 3'b000;
    assign _3861 = { _3860,
                     _271 };
    assign _3858 = { _3860,
                     _266 };
    assign _220 = 1'b0;
    assign _3452 = { _3860,
                     _276 };
    assign _3449 = { _3860,
                     _271 };
    assign _3446 = { _3860,
                     _266 };
    assign _3433 = { _3860,
                     _281 };
    assign _3430 = { _3860,
                     _276 };
    assign _3427 = { _3860,
                     _271 };
    assign _3414 = { _3860,
                     _286 };
    assign _3411 = { _3860,
                     _281 };
    assign _3408 = { _3860,
                     _276 };
    assign _3395 = { _3860,
                     _291 };
    assign _3392 = { _3860,
                     _286 };
    assign _3389 = { _3860,
                     _281 };
    assign _3376 = { _3860,
                     _296 };
    assign _3373 = { _3860,
                     _291 };
    assign _3370 = { _3860,
                     _286 };
    assign _3357 = { _3860,
                     _301 };
    assign _3354 = { _3860,
                     _296 };
    assign _3351 = { _3860,
                     _291 };
    assign _3338 = { _3860,
                     _306 };
    assign _3335 = { _3860,
                     _301 };
    assign _3332 = { _3860,
                     _296 };
    assign _3319 = { _3860,
                     _311 };
    assign _3316 = { _3860,
                     _306 };
    assign _3313 = { _3860,
                     _301 };
    assign _3300 = { _3860,
                     _311 };
    assign _3072 = { _3860,
                     _361 };
    assign _3069 = { _3860,
                     _356 };
    assign _3066 = { _3860,
                     _351 };
    assign _3063 = { _3860,
                     _311 };
    assign _3100 = { _3860,
                     _356 };
    assign _3097 = { _3860,
                     _351 };
    assign _3094 = { _3860,
                     _346 };
    assign _3091 = { _3860,
                     _306 };
    assign _3128 = { _3860,
                     _351 };
    assign _3125 = { _3860,
                     _346 };
    assign _3122 = { _3860,
                     _341 };
    assign _3119 = { _3860,
                     _301 };
    assign _3156 = { _3860,
                     _346 };
    assign _3153 = { _3860,
                     _341 };
    assign _3150 = { _3860,
                     _336 };
    assign _3147 = { _3860,
                     _296 };
    assign _3184 = { _3860,
                     _341 };
    assign _3181 = { _3860,
                     _336 };
    assign _3178 = { _3860,
                     _331 };
    assign _3175 = { _3860,
                     _291 };
    assign _3212 = { _3860,
                     _336 };
    assign _3209 = { _3860,
                     _331 };
    assign _3206 = { _3860,
                     _326 };
    assign _3203 = { _3860,
                     _286 };
    assign _3240 = { _3860,
                     _331 };
    assign _3237 = { _3860,
                     _326 };
    assign _3234 = { _3860,
                     _321 };
    assign _3231 = { _3860,
                     _281 };
    assign _3268 = { _3860,
                     _326 };
    assign _3265 = { _3860,
                     _321 };
    assign _3262 = { _3860,
                     _316 };
    assign _3259 = { _3860,
                     _276 };
    assign _3287 = { _3860,
                     _321 };
    assign _3025 = { _3860,
                     _371 };
    assign _3022 = { _3860,
                     _366 };
    assign _3006 = { _3860,
                     _376 };
    assign _3003 = { _3860,
                     _371 };
    assign _3000 = { _3860,
                     _366 };
    assign _2978 = { _3860,
                     _381 };
    assign _2975 = { _3860,
                     _376 };
    assign _2972 = { _3860,
                     _371 };
    assign _2950 = { _3860,
                     _386 };
    assign _2947 = { _3860,
                     _381 };
    assign _2944 = { _3860,
                     _376 };
    assign _2922 = { _3860,
                     _391 };
    assign _2919 = { _3860,
                     _386 };
    assign _2916 = { _3860,
                     _381 };
    assign _2894 = { _3860,
                     _396 };
    assign _2891 = { _3860,
                     _391 };
    assign _2888 = { _3860,
                     _386 };
    assign _2866 = { _3860,
                     _401 };
    assign _2863 = { _3860,
                     _396 };
    assign _2860 = { _3860,
                     _391 };
    assign _2838 = { _3860,
                     _406 };
    assign _2835 = { _3860,
                     _401 };
    assign _2832 = { _3860,
                     _396 };
    assign _2810 = { _3860,
                     _411 };
    assign _2807 = { _3860,
                     _406 };
    assign _2804 = { _3860,
                     _401 };
    assign _2801 = { _3860,
                     _361 };
    assign _2798 = { _3860,
                     _351 };
    assign _2782 = { _3860,
                     _411 };
    assign _2548 = { _3860,
                     _461 };
    assign _2545 = { _3860,
                     _456 };
    assign _2542 = { _3860,
                     _451 };
    assign _2539 = { _3860,
                     _411 };
    assign _2576 = { _3860,
                     _456 };
    assign _2573 = { _3860,
                     _451 };
    assign _2570 = { _3860,
                     _446 };
    assign _2567 = { _3860,
                     _406 };
    assign _2604 = { _3860,
                     _451 };
    assign _2601 = { _3860,
                     _446 };
    assign _2598 = { _3860,
                     _441 };
    assign _2595 = { _3860,
                     _401 };
    assign _2632 = { _3860,
                     _446 };
    assign _2629 = { _3860,
                     _441 };
    assign _2626 = { _3860,
                     _436 };
    assign _2623 = { _3860,
                     _396 };
    assign _2660 = { _3860,
                     _441 };
    assign _2657 = { _3860,
                     _436 };
    assign _2654 = { _3860,
                     _431 };
    assign _2651 = { _3860,
                     _391 };
    assign _2688 = { _3860,
                     _436 };
    assign _2685 = { _3860,
                     _431 };
    assign _2682 = { _3860,
                     _426 };
    assign _2679 = { _3860,
                     _386 };
    assign _2716 = { _3860,
                     _431 };
    assign _2713 = { _3860,
                     _426 };
    assign _2710 = { _3860,
                     _421 };
    assign _2707 = { _3860,
                     _381 };
    assign _2744 = { _3860,
                     _426 };
    assign _2741 = { _3860,
                     _421 };
    assign _2738 = { _3860,
                     _416 };
    assign _2735 = { _3860,
                     _376 };
    assign _2763 = { _3860,
                     _421 };
    assign _2501 = { _3860,
                     _471 };
    assign _2498 = { _3860,
                     _466 };
    assign _2482 = { _3860,
                     _476 };
    assign _2479 = { _3860,
                     _471 };
    assign _2476 = { _3860,
                     _466 };
    assign _2454 = { _3860,
                     _481 };
    assign _2451 = { _3860,
                     _476 };
    assign _2448 = { _3860,
                     _471 };
    assign _2426 = { _3860,
                     _486 };
    assign _2423 = { _3860,
                     _481 };
    assign _2420 = { _3860,
                     _476 };
    assign _2398 = { _3860,
                     _491 };
    assign _2395 = { _3860,
                     _486 };
    assign _2392 = { _3860,
                     _481 };
    assign _2370 = { _3860,
                     _496 };
    assign _2367 = { _3860,
                     _491 };
    assign _2364 = { _3860,
                     _486 };
    assign _2342 = { _3860,
                     _501 };
    assign _2339 = { _3860,
                     _496 };
    assign _2336 = { _3860,
                     _491 };
    assign _2314 = { _3860,
                     _506 };
    assign _2311 = { _3860,
                     _501 };
    assign _2308 = { _3860,
                     _496 };
    assign _2286 = { _3860,
                     _511 };
    assign _2283 = { _3860,
                     _506 };
    assign _2280 = { _3860,
                     _501 };
    assign _2277 = { _3860,
                     _461 };
    assign _2274 = { _3860,
                     _451 };
    assign _2258 = { _3860,
                     _511 };
    assign _2024 = { _3860,
                     _561 };
    assign _2021 = { _3860,
                     _556 };
    assign _2018 = { _3860,
                     _551 };
    assign _2015 = { _3860,
                     _511 };
    assign _2052 = { _3860,
                     _556 };
    assign _2049 = { _3860,
                     _551 };
    assign _2046 = { _3860,
                     _546 };
    assign _2043 = { _3860,
                     _506 };
    assign _2080 = { _3860,
                     _551 };
    assign _2077 = { _3860,
                     _546 };
    assign _2074 = { _3860,
                     _541 };
    assign _2071 = { _3860,
                     _501 };
    assign _2108 = { _3860,
                     _546 };
    assign _2105 = { _3860,
                     _541 };
    assign _2102 = { _3860,
                     _536 };
    assign _2099 = { _3860,
                     _496 };
    assign _2136 = { _3860,
                     _541 };
    assign _2133 = { _3860,
                     _536 };
    assign _2130 = { _3860,
                     _531 };
    assign _2127 = { _3860,
                     _491 };
    assign _2164 = { _3860,
                     _536 };
    assign _2161 = { _3860,
                     _531 };
    assign _2158 = { _3860,
                     _526 };
    assign _2155 = { _3860,
                     _486 };
    assign _2192 = { _3860,
                     _531 };
    assign _2189 = { _3860,
                     _526 };
    assign _2186 = { _3860,
                     _521 };
    assign _2183 = { _3860,
                     _481 };
    assign _2220 = { _3860,
                     _526 };
    assign _2217 = { _3860,
                     _521 };
    assign _2214 = { _3860,
                     _516 };
    assign _2211 = { _3860,
                     _476 };
    assign _2239 = { _3860,
                     _521 };
    assign _1977 = { _3860,
                     _571 };
    assign _1974 = { _3860,
                     _566 };
    assign _1958 = { _3860,
                     _576 };
    assign _1955 = { _3860,
                     _571 };
    assign _1952 = { _3860,
                     _566 };
    assign _1930 = { _3860,
                     _581 };
    assign _1927 = { _3860,
                     _576 };
    assign _1924 = { _3860,
                     _571 };
    assign _1902 = { _3860,
                     _586 };
    assign _1899 = { _3860,
                     _581 };
    assign _1896 = { _3860,
                     _576 };
    assign _1874 = { _3860,
                     _591 };
    assign _1871 = { _3860,
                     _586 };
    assign _1868 = { _3860,
                     _581 };
    assign _1846 = { _3860,
                     _596 };
    assign _1843 = { _3860,
                     _591 };
    assign _1840 = { _3860,
                     _586 };
    assign _1818 = { _3860,
                     _601 };
    assign _1815 = { _3860,
                     _596 };
    assign _1812 = { _3860,
                     _591 };
    assign _1790 = { _3860,
                     _606 };
    assign _1787 = { _3860,
                     _601 };
    assign _1784 = { _3860,
                     _596 };
    assign _1762 = { _3860,
                     _611 };
    assign _1759 = { _3860,
                     _606 };
    assign _1756 = { _3860,
                     _601 };
    assign _1753 = { _3860,
                     _561 };
    assign _1750 = { _3860,
                     _551 };
    assign _1734 = { _3860,
                     _611 };
    assign _1500 = { _3860,
                     _661 };
    assign _1497 = { _3860,
                     _656 };
    assign _1494 = { _3860,
                     _651 };
    assign _1491 = { _3860,
                     _611 };
    assign _1528 = { _3860,
                     _656 };
    assign _1525 = { _3860,
                     _651 };
    assign _1522 = { _3860,
                     _646 };
    assign _1519 = { _3860,
                     _606 };
    assign _1556 = { _3860,
                     _651 };
    assign _1553 = { _3860,
                     _646 };
    assign _1550 = { _3860,
                     _641 };
    assign _1547 = { _3860,
                     _601 };
    assign _1584 = { _3860,
                     _646 };
    assign _1581 = { _3860,
                     _641 };
    assign _1578 = { _3860,
                     _636 };
    assign _1575 = { _3860,
                     _596 };
    assign _1612 = { _3860,
                     _641 };
    assign _1609 = { _3860,
                     _636 };
    assign _1606 = { _3860,
                     _631 };
    assign _1603 = { _3860,
                     _591 };
    assign _1640 = { _3860,
                     _636 };
    assign _1637 = { _3860,
                     _631 };
    assign _1634 = { _3860,
                     _626 };
    assign _1631 = { _3860,
                     _586 };
    assign _1668 = { _3860,
                     _631 };
    assign _1665 = { _3860,
                     _626 };
    assign _1662 = { _3860,
                     _621 };
    assign _1659 = { _3860,
                     _581 };
    assign _1696 = { _3860,
                     _626 };
    assign _1693 = { _3860,
                     _621 };
    assign _1690 = { _3860,
                     _616 };
    assign _1687 = { _3860,
                     _576 };
    assign _1715 = { _3860,
                     _621 };
    assign _1453 = { _3860,
                     _671 };
    assign _1450 = { _3860,
                     _666 };
    assign _1434 = { _3860,
                     _676 };
    assign _1431 = { _3860,
                     _671 };
    assign _1428 = { _3860,
                     _666 };
    assign _1406 = { _3860,
                     _681 };
    assign _1403 = { _3860,
                     _676 };
    assign _1400 = { _3860,
                     _671 };
    assign _1378 = { _3860,
                     _686 };
    assign _1375 = { _3860,
                     _681 };
    assign _1372 = { _3860,
                     _676 };
    assign _1350 = { _3860,
                     _691 };
    assign _1347 = { _3860,
                     _686 };
    assign _1344 = { _3860,
                     _681 };
    assign _1322 = { _3860,
                     _696 };
    assign _1319 = { _3860,
                     _691 };
    assign _1316 = { _3860,
                     _686 };
    assign _1294 = { _3860,
                     _701 };
    assign _1291 = { _3860,
                     _696 };
    assign _1288 = { _3860,
                     _691 };
    assign _1266 = { _3860,
                     _706 };
    assign _1263 = { _3860,
                     _701 };
    assign _1260 = { _3860,
                     _696 };
    assign _1238 = { _3860,
                     _711 };
    assign _1235 = { _3860,
                     _706 };
    assign _1232 = { _3860,
                     _701 };
    assign _1229 = { _3860,
                     _661 };
    assign _1226 = { _3860,
                     _651 };
    assign _1210 = { _3860,
                     _711 };
    assign _1026 = { _3860,
                     _706 };
    assign _1023 = { _3860,
                     _661 };
    assign _1021 = { _3860,
                     _656 };
    assign _1024 = _1021 + _1023;
    assign _1027 = _1024 + _1026;
    assign _1029 = _1027 < _3863;
    assign _1030 = _711 & _1029;
    assign _3459 = ~ _1030;
    assign _3460 = _711 & _3459;
    assign _3461 = _213 ? _3460 : _711;
    assign _3462 = _210 ? _706 : _3461;
    assign _103 = _3462;
    always @(posedge _205) begin
        if (_203)
            _711 <= _220;
        else
            _711 <= _103;
    end
    assign _1045 = { _3860,
                     _711 };
    assign _1064 = { _3860,
                     _706 };
    assign _1083 = { _3860,
                     _701 };
    assign _1102 = { _3860,
                     _696 };
    assign _1121 = { _3860,
                     _691 };
    assign _1140 = { _3860,
                     _686 };
    assign _1159 = { _3860,
                     _681 };
    assign _1178 = { _3860,
                     _676 };
    assign _1191 = { _3860,
                     _671 };
    assign _1188 = { _3860,
                     _621 };
    assign _1186 = { _3860,
                     _616 };
    assign _1189 = _1186 + _1188;
    assign _1192 = _1189 + _1191;
    assign _1194 = _1192 < _3863;
    assign _1195 = _666 & _1194;
    assign _3463 = ~ _1195;
    assign _3464 = _666 & _3463;
    assign _3465 = _213 ? _3464 : _666;
    assign _3466 = _210 ? _661 : _3465;
    assign _104 = _3466;
    always @(posedge _205) begin
        if (_203)
            _666 <= _220;
        else
            _666 <= _104;
    end
    assign _1175 = { _3860,
                     _666 };
    assign _1172 = { _3860,
                     _626 };
    assign _1169 = { _3860,
                     _621 };
    assign _1167 = { _3860,
                     _616 };
    assign _1170 = _1167 + _1169;
    assign _1173 = _1170 + _1172;
    assign _1176 = _1173 + _1175;
    assign _1179 = _1176 + _1178;
    assign _1181 = _1179 < _3863;
    assign _1182 = _671 & _1181;
    assign _3467 = ~ _1182;
    assign _3468 = _671 & _3467;
    assign _3469 = _213 ? _3468 : _671;
    assign _3470 = _210 ? _666 : _3469;
    assign _105 = _3470;
    always @(posedge _205) begin
        if (_203)
            _671 <= _220;
        else
            _671 <= _105;
    end
    assign _1156 = { _3860,
                     _671 };
    assign _1153 = { _3860,
                     _631 };
    assign _1150 = { _3860,
                     _626 };
    assign _1148 = { _3860,
                     _621 };
    assign _1151 = _1148 + _1150;
    assign _1154 = _1151 + _1153;
    assign _1157 = _1154 + _1156;
    assign _1160 = _1157 + _1159;
    assign _1162 = _1160 < _3863;
    assign _1163 = _676 & _1162;
    assign _3471 = ~ _1163;
    assign _3472 = _676 & _3471;
    assign _3473 = _213 ? _3472 : _676;
    assign _3474 = _210 ? _671 : _3473;
    assign _106 = _3474;
    always @(posedge _205) begin
        if (_203)
            _676 <= _220;
        else
            _676 <= _106;
    end
    assign _1137 = { _3860,
                     _676 };
    assign _1134 = { _3860,
                     _636 };
    assign _1131 = { _3860,
                     _631 };
    assign _1129 = { _3860,
                     _626 };
    assign _1132 = _1129 + _1131;
    assign _1135 = _1132 + _1134;
    assign _1138 = _1135 + _1137;
    assign _1141 = _1138 + _1140;
    assign _1143 = _1141 < _3863;
    assign _1144 = _681 & _1143;
    assign _3475 = ~ _1144;
    assign _3476 = _681 & _3475;
    assign _3477 = _213 ? _3476 : _681;
    assign _3478 = _210 ? _676 : _3477;
    assign _107 = _3478;
    always @(posedge _205) begin
        if (_203)
            _681 <= _220;
        else
            _681 <= _107;
    end
    assign _1118 = { _3860,
                     _681 };
    assign _1115 = { _3860,
                     _641 };
    assign _1112 = { _3860,
                     _636 };
    assign _1110 = { _3860,
                     _631 };
    assign _1113 = _1110 + _1112;
    assign _1116 = _1113 + _1115;
    assign _1119 = _1116 + _1118;
    assign _1122 = _1119 + _1121;
    assign _1124 = _1122 < _3863;
    assign _1125 = _686 & _1124;
    assign _3479 = ~ _1125;
    assign _3480 = _686 & _3479;
    assign _3481 = _213 ? _3480 : _686;
    assign _3482 = _210 ? _681 : _3481;
    assign _108 = _3482;
    always @(posedge _205) begin
        if (_203)
            _686 <= _220;
        else
            _686 <= _108;
    end
    assign _1099 = { _3860,
                     _686 };
    assign _1096 = { _3860,
                     _646 };
    assign _1093 = { _3860,
                     _641 };
    assign _1091 = { _3860,
                     _636 };
    assign _1094 = _1091 + _1093;
    assign _1097 = _1094 + _1096;
    assign _1100 = _1097 + _1099;
    assign _1103 = _1100 + _1102;
    assign _1105 = _1103 < _3863;
    assign _1106 = _691 & _1105;
    assign _3483 = ~ _1106;
    assign _3484 = _691 & _3483;
    assign _3485 = _213 ? _3484 : _691;
    assign _3486 = _210 ? _686 : _3485;
    assign _109 = _3486;
    always @(posedge _205) begin
        if (_203)
            _691 <= _220;
        else
            _691 <= _109;
    end
    assign _1080 = { _3860,
                     _691 };
    assign _1077 = { _3860,
                     _651 };
    assign _1074 = { _3860,
                     _646 };
    assign _1072 = { _3860,
                     _641 };
    assign _1075 = _1072 + _1074;
    assign _1078 = _1075 + _1077;
    assign _1081 = _1078 + _1080;
    assign _1084 = _1081 + _1083;
    assign _1086 = _1084 < _3863;
    assign _1087 = _696 & _1086;
    assign _3487 = ~ _1087;
    assign _3488 = _696 & _3487;
    assign _3489 = _213 ? _3488 : _696;
    assign _3490 = _210 ? _691 : _3489;
    assign _110 = _3490;
    always @(posedge _205) begin
        if (_203)
            _696 <= _220;
        else
            _696 <= _110;
    end
    assign _1061 = { _3860,
                     _696 };
    assign _1058 = { _3860,
                     _656 };
    assign _1055 = { _3860,
                     _651 };
    assign _1053 = { _3860,
                     _646 };
    assign _1056 = _1053 + _1055;
    assign _1059 = _1056 + _1058;
    assign _1062 = _1059 + _1061;
    assign _1065 = _1062 + _1064;
    assign _1067 = _1065 < _3863;
    assign _1068 = _701 & _1067;
    assign _3491 = ~ _1068;
    assign _3492 = _701 & _3491;
    assign _3493 = _213 ? _3492 : _701;
    assign _3494 = _210 ? _696 : _3493;
    assign _111 = _3494;
    always @(posedge _205) begin
        if (_203)
            _701 <= _220;
        else
            _701 <= _111;
    end
    assign _1042 = { _3860,
                     _701 };
    assign _1039 = { _3860,
                     _661 };
    assign _1036 = { _3860,
                     _656 };
    assign _1034 = { _3860,
                     _651 };
    assign _1037 = _1034 + _1036;
    assign _1040 = _1037 + _1039;
    assign _1043 = _1040 + _1042;
    assign _1046 = _1043 + _1045;
    assign _1048 = _1046 < _3863;
    assign _1049 = _706 & _1048;
    assign _3495 = ~ _1049;
    assign _3496 = _706 & _3495;
    assign _3497 = _213 ? _3496 : _706;
    assign _3498 = _210 ? _701 : _3497;
    assign _112 = _3498;
    always @(posedge _205) begin
        if (_203)
            _706 <= _220;
        else
            _706 <= _112;
    end
    assign _1207 = { _3860,
                     _706 };
    assign _1204 = { _3860,
                     _656 };
    assign _1201 = { _3860,
                     _611 };
    assign _1199 = { _3860,
                     _606 };
    assign _1202 = _1199 + _1201;
    assign _1205 = _1202 + _1204;
    assign _1208 = _1205 + _1207;
    assign _1211 = _1208 + _1210;
    assign _1213 = _1211 < _3863;
    assign _1214 = _661 & _1213;
    assign _3499 = ~ _1214;
    assign _3500 = _661 & _3499;
    assign _3501 = _213 ? _3500 : _661;
    assign _3502 = _210 ? _656 : _3501;
    assign _113 = _3502;
    always @(posedge _205) begin
        if (_203)
            _661 <= _220;
        else
            _661 <= _113;
    end
    assign _1472 = { _3860,
                     _661 };
    assign _1469 = { _3860,
                     _656 };
    assign _1466 = { _3860,
                     _606 };
    assign _1463 = { _3860,
                     _561 };
    assign _1461 = { _3860,
                     _556 };
    assign _1464 = _1461 + _1463;
    assign _1467 = _1464 + _1466;
    assign _1470 = _1467 + _1469;
    assign _1473 = _1470 + _1472;
    assign _1475 = _1473 < _3863;
    assign _1476 = _611 & _1475;
    assign _3503 = ~ _1476;
    assign _3504 = _611 & _3503;
    assign _3505 = _213 ? _3504 : _611;
    assign _3506 = _210 ? _606 : _3505;
    assign _114 = _3506;
    always @(posedge _205) begin
        if (_203)
            _611 <= _220;
        else
            _611 <= _114;
    end
    assign _1223 = { _3860,
                     _611 };
    assign _1220 = { _3860,
                     _606 };
    assign _1218 = { _3860,
                     _601 };
    assign _1221 = _1218 + _1220;
    assign _1224 = _1221 + _1223;
    assign _1227 = _1224 + _1226;
    assign _1230 = _1227 + _1229;
    assign _1233 = _1230 + _1232;
    assign _1236 = _1233 + _1235;
    assign _1239 = _1236 + _1238;
    assign _1241 = _1239 < _3863;
    assign _1242 = _656 & _1241;
    assign _3507 = ~ _1242;
    assign _3508 = _656 & _3507;
    assign _3509 = _213 ? _3508 : _656;
    assign _3510 = _210 ? _651 : _3509;
    assign _115 = _3510;
    always @(posedge _205) begin
        if (_203)
            _656 <= _220;
        else
            _656 <= _115;
    end
    assign _1257 = { _3860,
                     _656 };
    assign _1254 = { _3860,
                     _646 };
    assign _1251 = { _3860,
                     _606 };
    assign _1248 = { _3860,
                     _601 };
    assign _1246 = { _3860,
                     _596 };
    assign _1249 = _1246 + _1248;
    assign _1252 = _1249 + _1251;
    assign _1255 = _1252 + _1254;
    assign _1258 = _1255 + _1257;
    assign _1261 = _1258 + _1260;
    assign _1264 = _1261 + _1263;
    assign _1267 = _1264 + _1266;
    assign _1269 = _1267 < _3863;
    assign _1270 = _651 & _1269;
    assign _3511 = ~ _1270;
    assign _3512 = _651 & _3511;
    assign _3513 = _213 ? _3512 : _651;
    assign _3514 = _210 ? _646 : _3513;
    assign _116 = _3514;
    always @(posedge _205) begin
        if (_203)
            _651 <= _220;
        else
            _651 <= _116;
    end
    assign _1285 = { _3860,
                     _651 };
    assign _1282 = { _3860,
                     _641 };
    assign _1279 = { _3860,
                     _601 };
    assign _1276 = { _3860,
                     _596 };
    assign _1274 = { _3860,
                     _591 };
    assign _1277 = _1274 + _1276;
    assign _1280 = _1277 + _1279;
    assign _1283 = _1280 + _1282;
    assign _1286 = _1283 + _1285;
    assign _1289 = _1286 + _1288;
    assign _1292 = _1289 + _1291;
    assign _1295 = _1292 + _1294;
    assign _1297 = _1295 < _3863;
    assign _1298 = _646 & _1297;
    assign _3515 = ~ _1298;
    assign _3516 = _646 & _3515;
    assign _3517 = _213 ? _3516 : _646;
    assign _3518 = _210 ? _641 : _3517;
    assign _117 = _3518;
    always @(posedge _205) begin
        if (_203)
            _646 <= _220;
        else
            _646 <= _117;
    end
    assign _1313 = { _3860,
                     _646 };
    assign _1310 = { _3860,
                     _636 };
    assign _1307 = { _3860,
                     _596 };
    assign _1304 = { _3860,
                     _591 };
    assign _1302 = { _3860,
                     _586 };
    assign _1305 = _1302 + _1304;
    assign _1308 = _1305 + _1307;
    assign _1311 = _1308 + _1310;
    assign _1314 = _1311 + _1313;
    assign _1317 = _1314 + _1316;
    assign _1320 = _1317 + _1319;
    assign _1323 = _1320 + _1322;
    assign _1325 = _1323 < _3863;
    assign _1326 = _641 & _1325;
    assign _3519 = ~ _1326;
    assign _3520 = _641 & _3519;
    assign _3521 = _213 ? _3520 : _641;
    assign _3522 = _210 ? _636 : _3521;
    assign _118 = _3522;
    always @(posedge _205) begin
        if (_203)
            _641 <= _220;
        else
            _641 <= _118;
    end
    assign _1341 = { _3860,
                     _641 };
    assign _1338 = { _3860,
                     _631 };
    assign _1335 = { _3860,
                     _591 };
    assign _1332 = { _3860,
                     _586 };
    assign _1330 = { _3860,
                     _581 };
    assign _1333 = _1330 + _1332;
    assign _1336 = _1333 + _1335;
    assign _1339 = _1336 + _1338;
    assign _1342 = _1339 + _1341;
    assign _1345 = _1342 + _1344;
    assign _1348 = _1345 + _1347;
    assign _1351 = _1348 + _1350;
    assign _1353 = _1351 < _3863;
    assign _1354 = _636 & _1353;
    assign _3523 = ~ _1354;
    assign _3524 = _636 & _3523;
    assign _3525 = _213 ? _3524 : _636;
    assign _3526 = _210 ? _631 : _3525;
    assign _119 = _3526;
    always @(posedge _205) begin
        if (_203)
            _636 <= _220;
        else
            _636 <= _119;
    end
    assign _1369 = { _3860,
                     _636 };
    assign _1366 = { _3860,
                     _626 };
    assign _1363 = { _3860,
                     _586 };
    assign _1360 = { _3860,
                     _581 };
    assign _1358 = { _3860,
                     _576 };
    assign _1361 = _1358 + _1360;
    assign _1364 = _1361 + _1363;
    assign _1367 = _1364 + _1366;
    assign _1370 = _1367 + _1369;
    assign _1373 = _1370 + _1372;
    assign _1376 = _1373 + _1375;
    assign _1379 = _1376 + _1378;
    assign _1381 = _1379 < _3863;
    assign _1382 = _631 & _1381;
    assign _3527 = ~ _1382;
    assign _3528 = _631 & _3527;
    assign _3529 = _213 ? _3528 : _631;
    assign _3530 = _210 ? _626 : _3529;
    assign _120 = _3530;
    always @(posedge _205) begin
        if (_203)
            _631 <= _220;
        else
            _631 <= _120;
    end
    assign _1397 = { _3860,
                     _631 };
    assign _1394 = { _3860,
                     _621 };
    assign _1391 = { _3860,
                     _581 };
    assign _1388 = { _3860,
                     _576 };
    assign _1386 = { _3860,
                     _571 };
    assign _1389 = _1386 + _1388;
    assign _1392 = _1389 + _1391;
    assign _1395 = _1392 + _1394;
    assign _1398 = _1395 + _1397;
    assign _1401 = _1398 + _1400;
    assign _1404 = _1401 + _1403;
    assign _1407 = _1404 + _1406;
    assign _1409 = _1407 < _3863;
    assign _1410 = _626 & _1409;
    assign _3531 = ~ _1410;
    assign _3532 = _626 & _3531;
    assign _3533 = _213 ? _3532 : _626;
    assign _3534 = _210 ? _621 : _3533;
    assign _121 = _3534;
    always @(posedge _205) begin
        if (_203)
            _626 <= _220;
        else
            _626 <= _121;
    end
    assign _1425 = { _3860,
                     _626 };
    assign _1422 = { _3860,
                     _616 };
    assign _1419 = { _3860,
                     _576 };
    assign _1416 = { _3860,
                     _571 };
    assign _1414 = { _3860,
                     _566 };
    assign _1417 = _1414 + _1416;
    assign _1420 = _1417 + _1419;
    assign _1423 = _1420 + _1422;
    assign _1426 = _1423 + _1425;
    assign _1429 = _1426 + _1428;
    assign _1432 = _1429 + _1431;
    assign _1435 = _1432 + _1434;
    assign _1437 = _1435 < _3863;
    assign _1438 = _621 & _1437;
    assign _3535 = ~ _1438;
    assign _3536 = _621 & _3535;
    assign _3537 = _213 ? _3536 : _621;
    assign _3538 = _210 ? _616 : _3537;
    assign _122 = _3538;
    always @(posedge _205) begin
        if (_203)
            _621 <= _220;
        else
            _621 <= _122;
    end
    assign _1447 = { _3860,
                     _621 };
    assign _1444 = { _3860,
                     _571 };
    assign _1442 = { _3860,
                     _566 };
    assign _1445 = _1442 + _1444;
    assign _1448 = _1445 + _1447;
    assign _1451 = _1448 + _1450;
    assign _1454 = _1451 + _1453;
    assign _1456 = _1454 < _3863;
    assign _1457 = _616 & _1456;
    assign _3539 = ~ _1457;
    assign _3540 = _616 & _3539;
    assign _3541 = _213 ? _3540 : _616;
    assign _3542 = _210 ? _611 : _3541;
    assign _123 = _3542;
    always @(posedge _205) begin
        if (_203)
            _616 <= _220;
        else
            _616 <= _123;
    end
    assign _1712 = { _3860,
                     _616 };
    assign _1709 = { _3860,
                     _571 };
    assign _1706 = { _3860,
                     _521 };
    assign _1704 = { _3860,
                     _516 };
    assign _1707 = _1704 + _1706;
    assign _1710 = _1707 + _1709;
    assign _1713 = _1710 + _1712;
    assign _1716 = _1713 + _1715;
    assign _1718 = _1716 < _3863;
    assign _1719 = _566 & _1718;
    assign _3543 = ~ _1719;
    assign _3544 = _566 & _3543;
    assign _3545 = _213 ? _3544 : _566;
    assign _3546 = _210 ? _561 : _3545;
    assign _124 = _3546;
    always @(posedge _205) begin
        if (_203)
            _566 <= _220;
        else
            _566 <= _124;
    end
    assign _1684 = { _3860,
                     _566 };
    assign _1681 = { _3860,
                     _526 };
    assign _1678 = { _3860,
                     _521 };
    assign _1676 = { _3860,
                     _516 };
    assign _1679 = _1676 + _1678;
    assign _1682 = _1679 + _1681;
    assign _1685 = _1682 + _1684;
    assign _1688 = _1685 + _1687;
    assign _1691 = _1688 + _1690;
    assign _1694 = _1691 + _1693;
    assign _1697 = _1694 + _1696;
    assign _1699 = _1697 < _3863;
    assign _1700 = _571 & _1699;
    assign _3547 = ~ _1700;
    assign _3548 = _571 & _3547;
    assign _3549 = _213 ? _3548 : _571;
    assign _3550 = _210 ? _566 : _3549;
    assign _125 = _3550;
    always @(posedge _205) begin
        if (_203)
            _571 <= _220;
        else
            _571 <= _125;
    end
    assign _1656 = { _3860,
                     _571 };
    assign _1653 = { _3860,
                     _531 };
    assign _1650 = { _3860,
                     _526 };
    assign _1648 = { _3860,
                     _521 };
    assign _1651 = _1648 + _1650;
    assign _1654 = _1651 + _1653;
    assign _1657 = _1654 + _1656;
    assign _1660 = _1657 + _1659;
    assign _1663 = _1660 + _1662;
    assign _1666 = _1663 + _1665;
    assign _1669 = _1666 + _1668;
    assign _1671 = _1669 < _3863;
    assign _1672 = _576 & _1671;
    assign _3551 = ~ _1672;
    assign _3552 = _576 & _3551;
    assign _3553 = _213 ? _3552 : _576;
    assign _3554 = _210 ? _571 : _3553;
    assign _126 = _3554;
    always @(posedge _205) begin
        if (_203)
            _576 <= _220;
        else
            _576 <= _126;
    end
    assign _1628 = { _3860,
                     _576 };
    assign _1625 = { _3860,
                     _536 };
    assign _1622 = { _3860,
                     _531 };
    assign _1620 = { _3860,
                     _526 };
    assign _1623 = _1620 + _1622;
    assign _1626 = _1623 + _1625;
    assign _1629 = _1626 + _1628;
    assign _1632 = _1629 + _1631;
    assign _1635 = _1632 + _1634;
    assign _1638 = _1635 + _1637;
    assign _1641 = _1638 + _1640;
    assign _1643 = _1641 < _3863;
    assign _1644 = _581 & _1643;
    assign _3555 = ~ _1644;
    assign _3556 = _581 & _3555;
    assign _3557 = _213 ? _3556 : _581;
    assign _3558 = _210 ? _576 : _3557;
    assign _127 = _3558;
    always @(posedge _205) begin
        if (_203)
            _581 <= _220;
        else
            _581 <= _127;
    end
    assign _1600 = { _3860,
                     _581 };
    assign _1597 = { _3860,
                     _541 };
    assign _1594 = { _3860,
                     _536 };
    assign _1592 = { _3860,
                     _531 };
    assign _1595 = _1592 + _1594;
    assign _1598 = _1595 + _1597;
    assign _1601 = _1598 + _1600;
    assign _1604 = _1601 + _1603;
    assign _1607 = _1604 + _1606;
    assign _1610 = _1607 + _1609;
    assign _1613 = _1610 + _1612;
    assign _1615 = _1613 < _3863;
    assign _1616 = _586 & _1615;
    assign _3559 = ~ _1616;
    assign _3560 = _586 & _3559;
    assign _3561 = _213 ? _3560 : _586;
    assign _3562 = _210 ? _581 : _3561;
    assign _128 = _3562;
    always @(posedge _205) begin
        if (_203)
            _586 <= _220;
        else
            _586 <= _128;
    end
    assign _1572 = { _3860,
                     _586 };
    assign _1569 = { _3860,
                     _546 };
    assign _1566 = { _3860,
                     _541 };
    assign _1564 = { _3860,
                     _536 };
    assign _1567 = _1564 + _1566;
    assign _1570 = _1567 + _1569;
    assign _1573 = _1570 + _1572;
    assign _1576 = _1573 + _1575;
    assign _1579 = _1576 + _1578;
    assign _1582 = _1579 + _1581;
    assign _1585 = _1582 + _1584;
    assign _1587 = _1585 < _3863;
    assign _1588 = _591 & _1587;
    assign _3563 = ~ _1588;
    assign _3564 = _591 & _3563;
    assign _3565 = _213 ? _3564 : _591;
    assign _3566 = _210 ? _586 : _3565;
    assign _129 = _3566;
    always @(posedge _205) begin
        if (_203)
            _591 <= _220;
        else
            _591 <= _129;
    end
    assign _1544 = { _3860,
                     _591 };
    assign _1541 = { _3860,
                     _551 };
    assign _1538 = { _3860,
                     _546 };
    assign _1536 = { _3860,
                     _541 };
    assign _1539 = _1536 + _1538;
    assign _1542 = _1539 + _1541;
    assign _1545 = _1542 + _1544;
    assign _1548 = _1545 + _1547;
    assign _1551 = _1548 + _1550;
    assign _1554 = _1551 + _1553;
    assign _1557 = _1554 + _1556;
    assign _1559 = _1557 < _3863;
    assign _1560 = _596 & _1559;
    assign _3567 = ~ _1560;
    assign _3568 = _596 & _3567;
    assign _3569 = _213 ? _3568 : _596;
    assign _3570 = _210 ? _591 : _3569;
    assign _130 = _3570;
    always @(posedge _205) begin
        if (_203)
            _596 <= _220;
        else
            _596 <= _130;
    end
    assign _1516 = { _3860,
                     _596 };
    assign _1513 = { _3860,
                     _556 };
    assign _1510 = { _3860,
                     _551 };
    assign _1508 = { _3860,
                     _546 };
    assign _1511 = _1508 + _1510;
    assign _1514 = _1511 + _1513;
    assign _1517 = _1514 + _1516;
    assign _1520 = _1517 + _1519;
    assign _1523 = _1520 + _1522;
    assign _1526 = _1523 + _1525;
    assign _1529 = _1526 + _1528;
    assign _1531 = _1529 < _3863;
    assign _1532 = _601 & _1531;
    assign _3571 = ~ _1532;
    assign _3572 = _601 & _3571;
    assign _3573 = _213 ? _3572 : _601;
    assign _3574 = _210 ? _596 : _3573;
    assign _131 = _3574;
    always @(posedge _205) begin
        if (_203)
            _601 <= _220;
        else
            _601 <= _131;
    end
    assign _1488 = { _3860,
                     _601 };
    assign _1485 = { _3860,
                     _561 };
    assign _1482 = { _3860,
                     _556 };
    assign _1480 = { _3860,
                     _551 };
    assign _1483 = _1480 + _1482;
    assign _1486 = _1483 + _1485;
    assign _1489 = _1486 + _1488;
    assign _1492 = _1489 + _1491;
    assign _1495 = _1492 + _1494;
    assign _1498 = _1495 + _1497;
    assign _1501 = _1498 + _1500;
    assign _1503 = _1501 < _3863;
    assign _1504 = _606 & _1503;
    assign _3575 = ~ _1504;
    assign _3576 = _606 & _3575;
    assign _3577 = _213 ? _3576 : _606;
    assign _3578 = _210 ? _601 : _3577;
    assign _132 = _3578;
    always @(posedge _205) begin
        if (_203)
            _606 <= _220;
        else
            _606 <= _132;
    end
    assign _1731 = { _3860,
                     _606 };
    assign _1728 = { _3860,
                     _556 };
    assign _1725 = { _3860,
                     _511 };
    assign _1723 = { _3860,
                     _506 };
    assign _1726 = _1723 + _1725;
    assign _1729 = _1726 + _1728;
    assign _1732 = _1729 + _1731;
    assign _1735 = _1732 + _1734;
    assign _1737 = _1735 < _3863;
    assign _1738 = _561 & _1737;
    assign _3579 = ~ _1738;
    assign _3580 = _561 & _3579;
    assign _3581 = _213 ? _3580 : _561;
    assign _3582 = _210 ? _556 : _3581;
    assign _133 = _3582;
    always @(posedge _205) begin
        if (_203)
            _561 <= _220;
        else
            _561 <= _133;
    end
    assign _1996 = { _3860,
                     _561 };
    assign _1993 = { _3860,
                     _556 };
    assign _1990 = { _3860,
                     _506 };
    assign _1987 = { _3860,
                     _461 };
    assign _1985 = { _3860,
                     _456 };
    assign _1988 = _1985 + _1987;
    assign _1991 = _1988 + _1990;
    assign _1994 = _1991 + _1993;
    assign _1997 = _1994 + _1996;
    assign _1999 = _1997 < _3863;
    assign _2000 = _511 & _1999;
    assign _3583 = ~ _2000;
    assign _3584 = _511 & _3583;
    assign _3585 = _213 ? _3584 : _511;
    assign _3586 = _210 ? _506 : _3585;
    assign _134 = _3586;
    always @(posedge _205) begin
        if (_203)
            _511 <= _220;
        else
            _511 <= _134;
    end
    assign _1747 = { _3860,
                     _511 };
    assign _1744 = { _3860,
                     _506 };
    assign _1742 = { _3860,
                     _501 };
    assign _1745 = _1742 + _1744;
    assign _1748 = _1745 + _1747;
    assign _1751 = _1748 + _1750;
    assign _1754 = _1751 + _1753;
    assign _1757 = _1754 + _1756;
    assign _1760 = _1757 + _1759;
    assign _1763 = _1760 + _1762;
    assign _1765 = _1763 < _3863;
    assign _1766 = _556 & _1765;
    assign _3587 = ~ _1766;
    assign _3588 = _556 & _3587;
    assign _3589 = _213 ? _3588 : _556;
    assign _3590 = _210 ? _551 : _3589;
    assign _135 = _3590;
    always @(posedge _205) begin
        if (_203)
            _556 <= _220;
        else
            _556 <= _135;
    end
    assign _1781 = { _3860,
                     _556 };
    assign _1778 = { _3860,
                     _546 };
    assign _1775 = { _3860,
                     _506 };
    assign _1772 = { _3860,
                     _501 };
    assign _1770 = { _3860,
                     _496 };
    assign _1773 = _1770 + _1772;
    assign _1776 = _1773 + _1775;
    assign _1779 = _1776 + _1778;
    assign _1782 = _1779 + _1781;
    assign _1785 = _1782 + _1784;
    assign _1788 = _1785 + _1787;
    assign _1791 = _1788 + _1790;
    assign _1793 = _1791 < _3863;
    assign _1794 = _551 & _1793;
    assign _3591 = ~ _1794;
    assign _3592 = _551 & _3591;
    assign _3593 = _213 ? _3592 : _551;
    assign _3594 = _210 ? _546 : _3593;
    assign _136 = _3594;
    always @(posedge _205) begin
        if (_203)
            _551 <= _220;
        else
            _551 <= _136;
    end
    assign _1809 = { _3860,
                     _551 };
    assign _1806 = { _3860,
                     _541 };
    assign _1803 = { _3860,
                     _501 };
    assign _1800 = { _3860,
                     _496 };
    assign _1798 = { _3860,
                     _491 };
    assign _1801 = _1798 + _1800;
    assign _1804 = _1801 + _1803;
    assign _1807 = _1804 + _1806;
    assign _1810 = _1807 + _1809;
    assign _1813 = _1810 + _1812;
    assign _1816 = _1813 + _1815;
    assign _1819 = _1816 + _1818;
    assign _1821 = _1819 < _3863;
    assign _1822 = _546 & _1821;
    assign _3595 = ~ _1822;
    assign _3596 = _546 & _3595;
    assign _3597 = _213 ? _3596 : _546;
    assign _3598 = _210 ? _541 : _3597;
    assign _137 = _3598;
    always @(posedge _205) begin
        if (_203)
            _546 <= _220;
        else
            _546 <= _137;
    end
    assign _1837 = { _3860,
                     _546 };
    assign _1834 = { _3860,
                     _536 };
    assign _1831 = { _3860,
                     _496 };
    assign _1828 = { _3860,
                     _491 };
    assign _1826 = { _3860,
                     _486 };
    assign _1829 = _1826 + _1828;
    assign _1832 = _1829 + _1831;
    assign _1835 = _1832 + _1834;
    assign _1838 = _1835 + _1837;
    assign _1841 = _1838 + _1840;
    assign _1844 = _1841 + _1843;
    assign _1847 = _1844 + _1846;
    assign _1849 = _1847 < _3863;
    assign _1850 = _541 & _1849;
    assign _3599 = ~ _1850;
    assign _3600 = _541 & _3599;
    assign _3601 = _213 ? _3600 : _541;
    assign _3602 = _210 ? _536 : _3601;
    assign _138 = _3602;
    always @(posedge _205) begin
        if (_203)
            _541 <= _220;
        else
            _541 <= _138;
    end
    assign _1865 = { _3860,
                     _541 };
    assign _1862 = { _3860,
                     _531 };
    assign _1859 = { _3860,
                     _491 };
    assign _1856 = { _3860,
                     _486 };
    assign _1854 = { _3860,
                     _481 };
    assign _1857 = _1854 + _1856;
    assign _1860 = _1857 + _1859;
    assign _1863 = _1860 + _1862;
    assign _1866 = _1863 + _1865;
    assign _1869 = _1866 + _1868;
    assign _1872 = _1869 + _1871;
    assign _1875 = _1872 + _1874;
    assign _1877 = _1875 < _3863;
    assign _1878 = _536 & _1877;
    assign _3603 = ~ _1878;
    assign _3604 = _536 & _3603;
    assign _3605 = _213 ? _3604 : _536;
    assign _3606 = _210 ? _531 : _3605;
    assign _139 = _3606;
    always @(posedge _205) begin
        if (_203)
            _536 <= _220;
        else
            _536 <= _139;
    end
    assign _1893 = { _3860,
                     _536 };
    assign _1890 = { _3860,
                     _526 };
    assign _1887 = { _3860,
                     _486 };
    assign _1884 = { _3860,
                     _481 };
    assign _1882 = { _3860,
                     _476 };
    assign _1885 = _1882 + _1884;
    assign _1888 = _1885 + _1887;
    assign _1891 = _1888 + _1890;
    assign _1894 = _1891 + _1893;
    assign _1897 = _1894 + _1896;
    assign _1900 = _1897 + _1899;
    assign _1903 = _1900 + _1902;
    assign _1905 = _1903 < _3863;
    assign _1906 = _531 & _1905;
    assign _3607 = ~ _1906;
    assign _3608 = _531 & _3607;
    assign _3609 = _213 ? _3608 : _531;
    assign _3610 = _210 ? _526 : _3609;
    assign _140 = _3610;
    always @(posedge _205) begin
        if (_203)
            _531 <= _220;
        else
            _531 <= _140;
    end
    assign _1921 = { _3860,
                     _531 };
    assign _1918 = { _3860,
                     _521 };
    assign _1915 = { _3860,
                     _481 };
    assign _1912 = { _3860,
                     _476 };
    assign _1910 = { _3860,
                     _471 };
    assign _1913 = _1910 + _1912;
    assign _1916 = _1913 + _1915;
    assign _1919 = _1916 + _1918;
    assign _1922 = _1919 + _1921;
    assign _1925 = _1922 + _1924;
    assign _1928 = _1925 + _1927;
    assign _1931 = _1928 + _1930;
    assign _1933 = _1931 < _3863;
    assign _1934 = _526 & _1933;
    assign _3611 = ~ _1934;
    assign _3612 = _526 & _3611;
    assign _3613 = _213 ? _3612 : _526;
    assign _3614 = _210 ? _521 : _3613;
    assign _141 = _3614;
    always @(posedge _205) begin
        if (_203)
            _526 <= _220;
        else
            _526 <= _141;
    end
    assign _1949 = { _3860,
                     _526 };
    assign _1946 = { _3860,
                     _516 };
    assign _1943 = { _3860,
                     _476 };
    assign _1940 = { _3860,
                     _471 };
    assign _1938 = { _3860,
                     _466 };
    assign _1941 = _1938 + _1940;
    assign _1944 = _1941 + _1943;
    assign _1947 = _1944 + _1946;
    assign _1950 = _1947 + _1949;
    assign _1953 = _1950 + _1952;
    assign _1956 = _1953 + _1955;
    assign _1959 = _1956 + _1958;
    assign _1961 = _1959 < _3863;
    assign _1962 = _521 & _1961;
    assign _3615 = ~ _1962;
    assign _3616 = _521 & _3615;
    assign _3617 = _213 ? _3616 : _521;
    assign _3618 = _210 ? _516 : _3617;
    assign _142 = _3618;
    always @(posedge _205) begin
        if (_203)
            _521 <= _220;
        else
            _521 <= _142;
    end
    assign _1971 = { _3860,
                     _521 };
    assign _1968 = { _3860,
                     _471 };
    assign _1966 = { _3860,
                     _466 };
    assign _1969 = _1966 + _1968;
    assign _1972 = _1969 + _1971;
    assign _1975 = _1972 + _1974;
    assign _1978 = _1975 + _1977;
    assign _1980 = _1978 < _3863;
    assign _1981 = _516 & _1980;
    assign _3619 = ~ _1981;
    assign _3620 = _516 & _3619;
    assign _3621 = _213 ? _3620 : _516;
    assign _3622 = _210 ? _511 : _3621;
    assign _143 = _3622;
    always @(posedge _205) begin
        if (_203)
            _516 <= _220;
        else
            _516 <= _143;
    end
    assign _2236 = { _3860,
                     _516 };
    assign _2233 = { _3860,
                     _471 };
    assign _2230 = { _3860,
                     _421 };
    assign _2228 = { _3860,
                     _416 };
    assign _2231 = _2228 + _2230;
    assign _2234 = _2231 + _2233;
    assign _2237 = _2234 + _2236;
    assign _2240 = _2237 + _2239;
    assign _2242 = _2240 < _3863;
    assign _2243 = _466 & _2242;
    assign _3623 = ~ _2243;
    assign _3624 = _466 & _3623;
    assign _3625 = _213 ? _3624 : _466;
    assign _3626 = _210 ? _461 : _3625;
    assign _144 = _3626;
    always @(posedge _205) begin
        if (_203)
            _466 <= _220;
        else
            _466 <= _144;
    end
    assign _2208 = { _3860,
                     _466 };
    assign _2205 = { _3860,
                     _426 };
    assign _2202 = { _3860,
                     _421 };
    assign _2200 = { _3860,
                     _416 };
    assign _2203 = _2200 + _2202;
    assign _2206 = _2203 + _2205;
    assign _2209 = _2206 + _2208;
    assign _2212 = _2209 + _2211;
    assign _2215 = _2212 + _2214;
    assign _2218 = _2215 + _2217;
    assign _2221 = _2218 + _2220;
    assign _2223 = _2221 < _3863;
    assign _2224 = _471 & _2223;
    assign _3627 = ~ _2224;
    assign _3628 = _471 & _3627;
    assign _3629 = _213 ? _3628 : _471;
    assign _3630 = _210 ? _466 : _3629;
    assign _145 = _3630;
    always @(posedge _205) begin
        if (_203)
            _471 <= _220;
        else
            _471 <= _145;
    end
    assign _2180 = { _3860,
                     _471 };
    assign _2177 = { _3860,
                     _431 };
    assign _2174 = { _3860,
                     _426 };
    assign _2172 = { _3860,
                     _421 };
    assign _2175 = _2172 + _2174;
    assign _2178 = _2175 + _2177;
    assign _2181 = _2178 + _2180;
    assign _2184 = _2181 + _2183;
    assign _2187 = _2184 + _2186;
    assign _2190 = _2187 + _2189;
    assign _2193 = _2190 + _2192;
    assign _2195 = _2193 < _3863;
    assign _2196 = _476 & _2195;
    assign _3631 = ~ _2196;
    assign _3632 = _476 & _3631;
    assign _3633 = _213 ? _3632 : _476;
    assign _3634 = _210 ? _471 : _3633;
    assign _146 = _3634;
    always @(posedge _205) begin
        if (_203)
            _476 <= _220;
        else
            _476 <= _146;
    end
    assign _2152 = { _3860,
                     _476 };
    assign _2149 = { _3860,
                     _436 };
    assign _2146 = { _3860,
                     _431 };
    assign _2144 = { _3860,
                     _426 };
    assign _2147 = _2144 + _2146;
    assign _2150 = _2147 + _2149;
    assign _2153 = _2150 + _2152;
    assign _2156 = _2153 + _2155;
    assign _2159 = _2156 + _2158;
    assign _2162 = _2159 + _2161;
    assign _2165 = _2162 + _2164;
    assign _2167 = _2165 < _3863;
    assign _2168 = _481 & _2167;
    assign _3635 = ~ _2168;
    assign _3636 = _481 & _3635;
    assign _3637 = _213 ? _3636 : _481;
    assign _3638 = _210 ? _476 : _3637;
    assign _147 = _3638;
    always @(posedge _205) begin
        if (_203)
            _481 <= _220;
        else
            _481 <= _147;
    end
    assign _2124 = { _3860,
                     _481 };
    assign _2121 = { _3860,
                     _441 };
    assign _2118 = { _3860,
                     _436 };
    assign _2116 = { _3860,
                     _431 };
    assign _2119 = _2116 + _2118;
    assign _2122 = _2119 + _2121;
    assign _2125 = _2122 + _2124;
    assign _2128 = _2125 + _2127;
    assign _2131 = _2128 + _2130;
    assign _2134 = _2131 + _2133;
    assign _2137 = _2134 + _2136;
    assign _2139 = _2137 < _3863;
    assign _2140 = _486 & _2139;
    assign _3639 = ~ _2140;
    assign _3640 = _486 & _3639;
    assign _3641 = _213 ? _3640 : _486;
    assign _3642 = _210 ? _481 : _3641;
    assign _148 = _3642;
    always @(posedge _205) begin
        if (_203)
            _486 <= _220;
        else
            _486 <= _148;
    end
    assign _2096 = { _3860,
                     _486 };
    assign _2093 = { _3860,
                     _446 };
    assign _2090 = { _3860,
                     _441 };
    assign _2088 = { _3860,
                     _436 };
    assign _2091 = _2088 + _2090;
    assign _2094 = _2091 + _2093;
    assign _2097 = _2094 + _2096;
    assign _2100 = _2097 + _2099;
    assign _2103 = _2100 + _2102;
    assign _2106 = _2103 + _2105;
    assign _2109 = _2106 + _2108;
    assign _2111 = _2109 < _3863;
    assign _2112 = _491 & _2111;
    assign _3643 = ~ _2112;
    assign _3644 = _491 & _3643;
    assign _3645 = _213 ? _3644 : _491;
    assign _3646 = _210 ? _486 : _3645;
    assign _149 = _3646;
    always @(posedge _205) begin
        if (_203)
            _491 <= _220;
        else
            _491 <= _149;
    end
    assign _2068 = { _3860,
                     _491 };
    assign _2065 = { _3860,
                     _451 };
    assign _2062 = { _3860,
                     _446 };
    assign _2060 = { _3860,
                     _441 };
    assign _2063 = _2060 + _2062;
    assign _2066 = _2063 + _2065;
    assign _2069 = _2066 + _2068;
    assign _2072 = _2069 + _2071;
    assign _2075 = _2072 + _2074;
    assign _2078 = _2075 + _2077;
    assign _2081 = _2078 + _2080;
    assign _2083 = _2081 < _3863;
    assign _2084 = _496 & _2083;
    assign _3647 = ~ _2084;
    assign _3648 = _496 & _3647;
    assign _3649 = _213 ? _3648 : _496;
    assign _3650 = _210 ? _491 : _3649;
    assign _150 = _3650;
    always @(posedge _205) begin
        if (_203)
            _496 <= _220;
        else
            _496 <= _150;
    end
    assign _2040 = { _3860,
                     _496 };
    assign _2037 = { _3860,
                     _456 };
    assign _2034 = { _3860,
                     _451 };
    assign _2032 = { _3860,
                     _446 };
    assign _2035 = _2032 + _2034;
    assign _2038 = _2035 + _2037;
    assign _2041 = _2038 + _2040;
    assign _2044 = _2041 + _2043;
    assign _2047 = _2044 + _2046;
    assign _2050 = _2047 + _2049;
    assign _2053 = _2050 + _2052;
    assign _2055 = _2053 < _3863;
    assign _2056 = _501 & _2055;
    assign _3651 = ~ _2056;
    assign _3652 = _501 & _3651;
    assign _3653 = _213 ? _3652 : _501;
    assign _3654 = _210 ? _496 : _3653;
    assign _151 = _3654;
    always @(posedge _205) begin
        if (_203)
            _501 <= _220;
        else
            _501 <= _151;
    end
    assign _2012 = { _3860,
                     _501 };
    assign _2009 = { _3860,
                     _461 };
    assign _2006 = { _3860,
                     _456 };
    assign _2004 = { _3860,
                     _451 };
    assign _2007 = _2004 + _2006;
    assign _2010 = _2007 + _2009;
    assign _2013 = _2010 + _2012;
    assign _2016 = _2013 + _2015;
    assign _2019 = _2016 + _2018;
    assign _2022 = _2019 + _2021;
    assign _2025 = _2022 + _2024;
    assign _2027 = _2025 < _3863;
    assign _2028 = _506 & _2027;
    assign _3655 = ~ _2028;
    assign _3656 = _506 & _3655;
    assign _3657 = _213 ? _3656 : _506;
    assign _3658 = _210 ? _501 : _3657;
    assign _152 = _3658;
    always @(posedge _205) begin
        if (_203)
            _506 <= _220;
        else
            _506 <= _152;
    end
    assign _2255 = { _3860,
                     _506 };
    assign _2252 = { _3860,
                     _456 };
    assign _2249 = { _3860,
                     _411 };
    assign _2247 = { _3860,
                     _406 };
    assign _2250 = _2247 + _2249;
    assign _2253 = _2250 + _2252;
    assign _2256 = _2253 + _2255;
    assign _2259 = _2256 + _2258;
    assign _2261 = _2259 < _3863;
    assign _2262 = _461 & _2261;
    assign _3659 = ~ _2262;
    assign _3660 = _461 & _3659;
    assign _3661 = _213 ? _3660 : _461;
    assign _3662 = _210 ? _456 : _3661;
    assign _153 = _3662;
    always @(posedge _205) begin
        if (_203)
            _461 <= _220;
        else
            _461 <= _153;
    end
    assign _2520 = { _3860,
                     _461 };
    assign _2517 = { _3860,
                     _456 };
    assign _2514 = { _3860,
                     _406 };
    assign _2511 = { _3860,
                     _361 };
    assign _2509 = { _3860,
                     _356 };
    assign _2512 = _2509 + _2511;
    assign _2515 = _2512 + _2514;
    assign _2518 = _2515 + _2517;
    assign _2521 = _2518 + _2520;
    assign _2523 = _2521 < _3863;
    assign _2524 = _411 & _2523;
    assign _3663 = ~ _2524;
    assign _3664 = _411 & _3663;
    assign _3665 = _213 ? _3664 : _411;
    assign _3666 = _210 ? _406 : _3665;
    assign _154 = _3666;
    always @(posedge _205) begin
        if (_203)
            _411 <= _220;
        else
            _411 <= _154;
    end
    assign _2271 = { _3860,
                     _411 };
    assign _2268 = { _3860,
                     _406 };
    assign _2266 = { _3860,
                     _401 };
    assign _2269 = _2266 + _2268;
    assign _2272 = _2269 + _2271;
    assign _2275 = _2272 + _2274;
    assign _2278 = _2275 + _2277;
    assign _2281 = _2278 + _2280;
    assign _2284 = _2281 + _2283;
    assign _2287 = _2284 + _2286;
    assign _2289 = _2287 < _3863;
    assign _2290 = _456 & _2289;
    assign _3667 = ~ _2290;
    assign _3668 = _456 & _3667;
    assign _3669 = _213 ? _3668 : _456;
    assign _3670 = _210 ? _451 : _3669;
    assign _155 = _3670;
    always @(posedge _205) begin
        if (_203)
            _456 <= _220;
        else
            _456 <= _155;
    end
    assign _2305 = { _3860,
                     _456 };
    assign _2302 = { _3860,
                     _446 };
    assign _2299 = { _3860,
                     _406 };
    assign _2296 = { _3860,
                     _401 };
    assign _2294 = { _3860,
                     _396 };
    assign _2297 = _2294 + _2296;
    assign _2300 = _2297 + _2299;
    assign _2303 = _2300 + _2302;
    assign _2306 = _2303 + _2305;
    assign _2309 = _2306 + _2308;
    assign _2312 = _2309 + _2311;
    assign _2315 = _2312 + _2314;
    assign _2317 = _2315 < _3863;
    assign _2318 = _451 & _2317;
    assign _3671 = ~ _2318;
    assign _3672 = _451 & _3671;
    assign _3673 = _213 ? _3672 : _451;
    assign _3674 = _210 ? _446 : _3673;
    assign _156 = _3674;
    always @(posedge _205) begin
        if (_203)
            _451 <= _220;
        else
            _451 <= _156;
    end
    assign _2333 = { _3860,
                     _451 };
    assign _2330 = { _3860,
                     _441 };
    assign _2327 = { _3860,
                     _401 };
    assign _2324 = { _3860,
                     _396 };
    assign _2322 = { _3860,
                     _391 };
    assign _2325 = _2322 + _2324;
    assign _2328 = _2325 + _2327;
    assign _2331 = _2328 + _2330;
    assign _2334 = _2331 + _2333;
    assign _2337 = _2334 + _2336;
    assign _2340 = _2337 + _2339;
    assign _2343 = _2340 + _2342;
    assign _2345 = _2343 < _3863;
    assign _2346 = _446 & _2345;
    assign _3675 = ~ _2346;
    assign _3676 = _446 & _3675;
    assign _3677 = _213 ? _3676 : _446;
    assign _3678 = _210 ? _441 : _3677;
    assign _157 = _3678;
    always @(posedge _205) begin
        if (_203)
            _446 <= _220;
        else
            _446 <= _157;
    end
    assign _2361 = { _3860,
                     _446 };
    assign _2358 = { _3860,
                     _436 };
    assign _2355 = { _3860,
                     _396 };
    assign _2352 = { _3860,
                     _391 };
    assign _2350 = { _3860,
                     _386 };
    assign _2353 = _2350 + _2352;
    assign _2356 = _2353 + _2355;
    assign _2359 = _2356 + _2358;
    assign _2362 = _2359 + _2361;
    assign _2365 = _2362 + _2364;
    assign _2368 = _2365 + _2367;
    assign _2371 = _2368 + _2370;
    assign _2373 = _2371 < _3863;
    assign _2374 = _441 & _2373;
    assign _3679 = ~ _2374;
    assign _3680 = _441 & _3679;
    assign _3681 = _213 ? _3680 : _441;
    assign _3682 = _210 ? _436 : _3681;
    assign _158 = _3682;
    always @(posedge _205) begin
        if (_203)
            _441 <= _220;
        else
            _441 <= _158;
    end
    assign _2389 = { _3860,
                     _441 };
    assign _2386 = { _3860,
                     _431 };
    assign _2383 = { _3860,
                     _391 };
    assign _2380 = { _3860,
                     _386 };
    assign _2378 = { _3860,
                     _381 };
    assign _2381 = _2378 + _2380;
    assign _2384 = _2381 + _2383;
    assign _2387 = _2384 + _2386;
    assign _2390 = _2387 + _2389;
    assign _2393 = _2390 + _2392;
    assign _2396 = _2393 + _2395;
    assign _2399 = _2396 + _2398;
    assign _2401 = _2399 < _3863;
    assign _2402 = _436 & _2401;
    assign _3683 = ~ _2402;
    assign _3684 = _436 & _3683;
    assign _3685 = _213 ? _3684 : _436;
    assign _3686 = _210 ? _431 : _3685;
    assign _159 = _3686;
    always @(posedge _205) begin
        if (_203)
            _436 <= _220;
        else
            _436 <= _159;
    end
    assign _2417 = { _3860,
                     _436 };
    assign _2414 = { _3860,
                     _426 };
    assign _2411 = { _3860,
                     _386 };
    assign _2408 = { _3860,
                     _381 };
    assign _2406 = { _3860,
                     _376 };
    assign _2409 = _2406 + _2408;
    assign _2412 = _2409 + _2411;
    assign _2415 = _2412 + _2414;
    assign _2418 = _2415 + _2417;
    assign _2421 = _2418 + _2420;
    assign _2424 = _2421 + _2423;
    assign _2427 = _2424 + _2426;
    assign _2429 = _2427 < _3863;
    assign _2430 = _431 & _2429;
    assign _3687 = ~ _2430;
    assign _3688 = _431 & _3687;
    assign _3689 = _213 ? _3688 : _431;
    assign _3690 = _210 ? _426 : _3689;
    assign _160 = _3690;
    always @(posedge _205) begin
        if (_203)
            _431 <= _220;
        else
            _431 <= _160;
    end
    assign _2445 = { _3860,
                     _431 };
    assign _2442 = { _3860,
                     _421 };
    assign _2439 = { _3860,
                     _381 };
    assign _2436 = { _3860,
                     _376 };
    assign _2434 = { _3860,
                     _371 };
    assign _2437 = _2434 + _2436;
    assign _2440 = _2437 + _2439;
    assign _2443 = _2440 + _2442;
    assign _2446 = _2443 + _2445;
    assign _2449 = _2446 + _2448;
    assign _2452 = _2449 + _2451;
    assign _2455 = _2452 + _2454;
    assign _2457 = _2455 < _3863;
    assign _2458 = _426 & _2457;
    assign _3691 = ~ _2458;
    assign _3692 = _426 & _3691;
    assign _3693 = _213 ? _3692 : _426;
    assign _3694 = _210 ? _421 : _3693;
    assign _161 = _3694;
    always @(posedge _205) begin
        if (_203)
            _426 <= _220;
        else
            _426 <= _161;
    end
    assign _2473 = { _3860,
                     _426 };
    assign _2470 = { _3860,
                     _416 };
    assign _2467 = { _3860,
                     _376 };
    assign _2464 = { _3860,
                     _371 };
    assign _2462 = { _3860,
                     _366 };
    assign _2465 = _2462 + _2464;
    assign _2468 = _2465 + _2467;
    assign _2471 = _2468 + _2470;
    assign _2474 = _2471 + _2473;
    assign _2477 = _2474 + _2476;
    assign _2480 = _2477 + _2479;
    assign _2483 = _2480 + _2482;
    assign _2485 = _2483 < _3863;
    assign _2486 = _421 & _2485;
    assign _3695 = ~ _2486;
    assign _3696 = _421 & _3695;
    assign _3697 = _213 ? _3696 : _421;
    assign _3698 = _210 ? _416 : _3697;
    assign _162 = _3698;
    always @(posedge _205) begin
        if (_203)
            _421 <= _220;
        else
            _421 <= _162;
    end
    assign _2495 = { _3860,
                     _421 };
    assign _2492 = { _3860,
                     _371 };
    assign _2490 = { _3860,
                     _366 };
    assign _2493 = _2490 + _2492;
    assign _2496 = _2493 + _2495;
    assign _2499 = _2496 + _2498;
    assign _2502 = _2499 + _2501;
    assign _2504 = _2502 < _3863;
    assign _2505 = _416 & _2504;
    assign _3699 = ~ _2505;
    assign _3700 = _416 & _3699;
    assign _3701 = _213 ? _3700 : _416;
    assign _3702 = _210 ? _411 : _3701;
    assign _163 = _3702;
    always @(posedge _205) begin
        if (_203)
            _416 <= _220;
        else
            _416 <= _163;
    end
    assign _2760 = { _3860,
                     _416 };
    assign _2757 = { _3860,
                     _371 };
    assign _2754 = { _3860,
                     _321 };
    assign _2752 = { _3860,
                     _316 };
    assign _2755 = _2752 + _2754;
    assign _2758 = _2755 + _2757;
    assign _2761 = _2758 + _2760;
    assign _2764 = _2761 + _2763;
    assign _2766 = _2764 < _3863;
    assign _2767 = _366 & _2766;
    assign _3703 = ~ _2767;
    assign _3704 = _366 & _3703;
    assign _3705 = _213 ? _3704 : _366;
    assign _3706 = _210 ? _361 : _3705;
    assign _164 = _3706;
    always @(posedge _205) begin
        if (_203)
            _366 <= _220;
        else
            _366 <= _164;
    end
    assign _2732 = { _3860,
                     _366 };
    assign _2729 = { _3860,
                     _326 };
    assign _2726 = { _3860,
                     _321 };
    assign _2724 = { _3860,
                     _316 };
    assign _2727 = _2724 + _2726;
    assign _2730 = _2727 + _2729;
    assign _2733 = _2730 + _2732;
    assign _2736 = _2733 + _2735;
    assign _2739 = _2736 + _2738;
    assign _2742 = _2739 + _2741;
    assign _2745 = _2742 + _2744;
    assign _2747 = _2745 < _3863;
    assign _2748 = _371 & _2747;
    assign _3707 = ~ _2748;
    assign _3708 = _371 & _3707;
    assign _3709 = _213 ? _3708 : _371;
    assign _3710 = _210 ? _366 : _3709;
    assign _165 = _3710;
    always @(posedge _205) begin
        if (_203)
            _371 <= _220;
        else
            _371 <= _165;
    end
    assign _2704 = { _3860,
                     _371 };
    assign _2701 = { _3860,
                     _331 };
    assign _2698 = { _3860,
                     _326 };
    assign _2696 = { _3860,
                     _321 };
    assign _2699 = _2696 + _2698;
    assign _2702 = _2699 + _2701;
    assign _2705 = _2702 + _2704;
    assign _2708 = _2705 + _2707;
    assign _2711 = _2708 + _2710;
    assign _2714 = _2711 + _2713;
    assign _2717 = _2714 + _2716;
    assign _2719 = _2717 < _3863;
    assign _2720 = _376 & _2719;
    assign _3711 = ~ _2720;
    assign _3712 = _376 & _3711;
    assign _3713 = _213 ? _3712 : _376;
    assign _3714 = _210 ? _371 : _3713;
    assign _166 = _3714;
    always @(posedge _205) begin
        if (_203)
            _376 <= _220;
        else
            _376 <= _166;
    end
    assign _2676 = { _3860,
                     _376 };
    assign _2673 = { _3860,
                     _336 };
    assign _2670 = { _3860,
                     _331 };
    assign _2668 = { _3860,
                     _326 };
    assign _2671 = _2668 + _2670;
    assign _2674 = _2671 + _2673;
    assign _2677 = _2674 + _2676;
    assign _2680 = _2677 + _2679;
    assign _2683 = _2680 + _2682;
    assign _2686 = _2683 + _2685;
    assign _2689 = _2686 + _2688;
    assign _2691 = _2689 < _3863;
    assign _2692 = _381 & _2691;
    assign _3715 = ~ _2692;
    assign _3716 = _381 & _3715;
    assign _3717 = _213 ? _3716 : _381;
    assign _3718 = _210 ? _376 : _3717;
    assign _167 = _3718;
    always @(posedge _205) begin
        if (_203)
            _381 <= _220;
        else
            _381 <= _167;
    end
    assign _2648 = { _3860,
                     _381 };
    assign _2645 = { _3860,
                     _341 };
    assign _2642 = { _3860,
                     _336 };
    assign _2640 = { _3860,
                     _331 };
    assign _2643 = _2640 + _2642;
    assign _2646 = _2643 + _2645;
    assign _2649 = _2646 + _2648;
    assign _2652 = _2649 + _2651;
    assign _2655 = _2652 + _2654;
    assign _2658 = _2655 + _2657;
    assign _2661 = _2658 + _2660;
    assign _2663 = _2661 < _3863;
    assign _2664 = _386 & _2663;
    assign _3719 = ~ _2664;
    assign _3720 = _386 & _3719;
    assign _3721 = _213 ? _3720 : _386;
    assign _3722 = _210 ? _381 : _3721;
    assign _168 = _3722;
    always @(posedge _205) begin
        if (_203)
            _386 <= _220;
        else
            _386 <= _168;
    end
    assign _2620 = { _3860,
                     _386 };
    assign _2617 = { _3860,
                     _346 };
    assign _2614 = { _3860,
                     _341 };
    assign _2612 = { _3860,
                     _336 };
    assign _2615 = _2612 + _2614;
    assign _2618 = _2615 + _2617;
    assign _2621 = _2618 + _2620;
    assign _2624 = _2621 + _2623;
    assign _2627 = _2624 + _2626;
    assign _2630 = _2627 + _2629;
    assign _2633 = _2630 + _2632;
    assign _2635 = _2633 < _3863;
    assign _2636 = _391 & _2635;
    assign _3723 = ~ _2636;
    assign _3724 = _391 & _3723;
    assign _3725 = _213 ? _3724 : _391;
    assign _3726 = _210 ? _386 : _3725;
    assign _169 = _3726;
    always @(posedge _205) begin
        if (_203)
            _391 <= _220;
        else
            _391 <= _169;
    end
    assign _2592 = { _3860,
                     _391 };
    assign _2589 = { _3860,
                     _351 };
    assign _2586 = { _3860,
                     _346 };
    assign _2584 = { _3860,
                     _341 };
    assign _2587 = _2584 + _2586;
    assign _2590 = _2587 + _2589;
    assign _2593 = _2590 + _2592;
    assign _2596 = _2593 + _2595;
    assign _2599 = _2596 + _2598;
    assign _2602 = _2599 + _2601;
    assign _2605 = _2602 + _2604;
    assign _2607 = _2605 < _3863;
    assign _2608 = _396 & _2607;
    assign _3727 = ~ _2608;
    assign _3728 = _396 & _3727;
    assign _3729 = _213 ? _3728 : _396;
    assign _3730 = _210 ? _391 : _3729;
    assign _170 = _3730;
    always @(posedge _205) begin
        if (_203)
            _396 <= _220;
        else
            _396 <= _170;
    end
    assign _2564 = { _3860,
                     _396 };
    assign _2561 = { _3860,
                     _356 };
    assign _2558 = { _3860,
                     _351 };
    assign _2556 = { _3860,
                     _346 };
    assign _2559 = _2556 + _2558;
    assign _2562 = _2559 + _2561;
    assign _2565 = _2562 + _2564;
    assign _2568 = _2565 + _2567;
    assign _2571 = _2568 + _2570;
    assign _2574 = _2571 + _2573;
    assign _2577 = _2574 + _2576;
    assign _2579 = _2577 < _3863;
    assign _2580 = _401 & _2579;
    assign _3731 = ~ _2580;
    assign _3732 = _401 & _3731;
    assign _3733 = _213 ? _3732 : _401;
    assign _3734 = _210 ? _396 : _3733;
    assign _171 = _3734;
    always @(posedge _205) begin
        if (_203)
            _401 <= _220;
        else
            _401 <= _171;
    end
    assign _2536 = { _3860,
                     _401 };
    assign _2533 = { _3860,
                     _361 };
    assign _2530 = { _3860,
                     _356 };
    assign _2528 = { _3860,
                     _351 };
    assign _2531 = _2528 + _2530;
    assign _2534 = _2531 + _2533;
    assign _2537 = _2534 + _2536;
    assign _2540 = _2537 + _2539;
    assign _2543 = _2540 + _2542;
    assign _2546 = _2543 + _2545;
    assign _2549 = _2546 + _2548;
    assign _2551 = _2549 < _3863;
    assign _2552 = _406 & _2551;
    assign _3735 = ~ _2552;
    assign _3736 = _406 & _3735;
    assign _3737 = _213 ? _3736 : _406;
    assign _3738 = _210 ? _401 : _3737;
    assign _172 = _3738;
    always @(posedge _205) begin
        if (_203)
            _406 <= _220;
        else
            _406 <= _172;
    end
    assign _2779 = { _3860,
                     _406 };
    assign _2776 = { _3860,
                     _356 };
    assign _2773 = { _3860,
                     _311 };
    assign _2771 = { _3860,
                     _306 };
    assign _2774 = _2771 + _2773;
    assign _2777 = _2774 + _2776;
    assign _2780 = _2777 + _2779;
    assign _2783 = _2780 + _2782;
    assign _2785 = _2783 < _3863;
    assign _2786 = _361 & _2785;
    assign _3739 = ~ _2786;
    assign _3740 = _361 & _3739;
    assign _3741 = _213 ? _3740 : _361;
    assign _3742 = _210 ? _356 : _3741;
    assign _173 = _3742;
    always @(posedge _205) begin
        if (_203)
            _361 <= _220;
        else
            _361 <= _173;
    end
    assign _3044 = { _3860,
                     _361 };
    assign _3041 = { _3860,
                     _356 };
    assign _3038 = { _3860,
                     _306 };
    assign _3035 = { _3860,
                     _261 };
    assign _3033 = { _3860,
                     _256 };
    assign _3036 = _3033 + _3035;
    assign _3039 = _3036 + _3038;
    assign _3042 = _3039 + _3041;
    assign _3045 = _3042 + _3044;
    assign _3047 = _3045 < _3863;
    assign _3048 = _311 & _3047;
    assign _3743 = ~ _3048;
    assign _3744 = _311 & _3743;
    assign _3745 = _213 ? _3744 : _311;
    assign _3746 = _210 ? _306 : _3745;
    assign _174 = _3746;
    always @(posedge _205) begin
        if (_203)
            _311 <= _220;
        else
            _311 <= _174;
    end
    assign _2795 = { _3860,
                     _311 };
    assign _2792 = { _3860,
                     _306 };
    assign _2790 = { _3860,
                     _301 };
    assign _2793 = _2790 + _2792;
    assign _2796 = _2793 + _2795;
    assign _2799 = _2796 + _2798;
    assign _2802 = _2799 + _2801;
    assign _2805 = _2802 + _2804;
    assign _2808 = _2805 + _2807;
    assign _2811 = _2808 + _2810;
    assign _2813 = _2811 < _3863;
    assign _2814 = _356 & _2813;
    assign _3747 = ~ _2814;
    assign _3748 = _356 & _3747;
    assign _3749 = _213 ? _3748 : _356;
    assign _3750 = _210 ? _351 : _3749;
    assign _175 = _3750;
    always @(posedge _205) begin
        if (_203)
            _356 <= _220;
        else
            _356 <= _175;
    end
    assign _2829 = { _3860,
                     _356 };
    assign _2826 = { _3860,
                     _346 };
    assign _2823 = { _3860,
                     _306 };
    assign _2820 = { _3860,
                     _301 };
    assign _2818 = { _3860,
                     _296 };
    assign _2821 = _2818 + _2820;
    assign _2824 = _2821 + _2823;
    assign _2827 = _2824 + _2826;
    assign _2830 = _2827 + _2829;
    assign _2833 = _2830 + _2832;
    assign _2836 = _2833 + _2835;
    assign _2839 = _2836 + _2838;
    assign _2841 = _2839 < _3863;
    assign _2842 = _351 & _2841;
    assign _3751 = ~ _2842;
    assign _3752 = _351 & _3751;
    assign _3753 = _213 ? _3752 : _351;
    assign _3754 = _210 ? _346 : _3753;
    assign _176 = _3754;
    always @(posedge _205) begin
        if (_203)
            _351 <= _220;
        else
            _351 <= _176;
    end
    assign _2857 = { _3860,
                     _351 };
    assign _2854 = { _3860,
                     _341 };
    assign _2851 = { _3860,
                     _301 };
    assign _2848 = { _3860,
                     _296 };
    assign _2846 = { _3860,
                     _291 };
    assign _2849 = _2846 + _2848;
    assign _2852 = _2849 + _2851;
    assign _2855 = _2852 + _2854;
    assign _2858 = _2855 + _2857;
    assign _2861 = _2858 + _2860;
    assign _2864 = _2861 + _2863;
    assign _2867 = _2864 + _2866;
    assign _2869 = _2867 < _3863;
    assign _2870 = _346 & _2869;
    assign _3755 = ~ _2870;
    assign _3756 = _346 & _3755;
    assign _3757 = _213 ? _3756 : _346;
    assign _3758 = _210 ? _341 : _3757;
    assign _177 = _3758;
    always @(posedge _205) begin
        if (_203)
            _346 <= _220;
        else
            _346 <= _177;
    end
    assign _2885 = { _3860,
                     _346 };
    assign _2882 = { _3860,
                     _336 };
    assign _2879 = { _3860,
                     _296 };
    assign _2876 = { _3860,
                     _291 };
    assign _2874 = { _3860,
                     _286 };
    assign _2877 = _2874 + _2876;
    assign _2880 = _2877 + _2879;
    assign _2883 = _2880 + _2882;
    assign _2886 = _2883 + _2885;
    assign _2889 = _2886 + _2888;
    assign _2892 = _2889 + _2891;
    assign _2895 = _2892 + _2894;
    assign _2897 = _2895 < _3863;
    assign _2898 = _341 & _2897;
    assign _3759 = ~ _2898;
    assign _3760 = _341 & _3759;
    assign _3761 = _213 ? _3760 : _341;
    assign _3762 = _210 ? _336 : _3761;
    assign _178 = _3762;
    always @(posedge _205) begin
        if (_203)
            _341 <= _220;
        else
            _341 <= _178;
    end
    assign _2913 = { _3860,
                     _341 };
    assign _2910 = { _3860,
                     _331 };
    assign _2907 = { _3860,
                     _291 };
    assign _2904 = { _3860,
                     _286 };
    assign _2902 = { _3860,
                     _281 };
    assign _2905 = _2902 + _2904;
    assign _2908 = _2905 + _2907;
    assign _2911 = _2908 + _2910;
    assign _2914 = _2911 + _2913;
    assign _2917 = _2914 + _2916;
    assign _2920 = _2917 + _2919;
    assign _2923 = _2920 + _2922;
    assign _2925 = _2923 < _3863;
    assign _2926 = _336 & _2925;
    assign _3763 = ~ _2926;
    assign _3764 = _336 & _3763;
    assign _3765 = _213 ? _3764 : _336;
    assign _3766 = _210 ? _331 : _3765;
    assign _179 = _3766;
    always @(posedge _205) begin
        if (_203)
            _336 <= _220;
        else
            _336 <= _179;
    end
    assign _2941 = { _3860,
                     _336 };
    assign _2938 = { _3860,
                     _326 };
    assign _2935 = { _3860,
                     _286 };
    assign _2932 = { _3860,
                     _281 };
    assign _2930 = { _3860,
                     _276 };
    assign _2933 = _2930 + _2932;
    assign _2936 = _2933 + _2935;
    assign _2939 = _2936 + _2938;
    assign _2942 = _2939 + _2941;
    assign _2945 = _2942 + _2944;
    assign _2948 = _2945 + _2947;
    assign _2951 = _2948 + _2950;
    assign _2953 = _2951 < _3863;
    assign _2954 = _331 & _2953;
    assign _3767 = ~ _2954;
    assign _3768 = _331 & _3767;
    assign _3769 = _213 ? _3768 : _331;
    assign _3770 = _210 ? _326 : _3769;
    assign _180 = _3770;
    always @(posedge _205) begin
        if (_203)
            _331 <= _220;
        else
            _331 <= _180;
    end
    assign _2969 = { _3860,
                     _331 };
    assign _2966 = { _3860,
                     _321 };
    assign _2963 = { _3860,
                     _281 };
    assign _2960 = { _3860,
                     _276 };
    assign _2958 = { _3860,
                     _271 };
    assign _2961 = _2958 + _2960;
    assign _2964 = _2961 + _2963;
    assign _2967 = _2964 + _2966;
    assign _2970 = _2967 + _2969;
    assign _2973 = _2970 + _2972;
    assign _2976 = _2973 + _2975;
    assign _2979 = _2976 + _2978;
    assign _2981 = _2979 < _3863;
    assign _2982 = _326 & _2981;
    assign _3771 = ~ _2982;
    assign _3772 = _326 & _3771;
    assign _3773 = _213 ? _3772 : _326;
    assign _3774 = _210 ? _321 : _3773;
    assign _181 = _3774;
    always @(posedge _205) begin
        if (_203)
            _326 <= _220;
        else
            _326 <= _181;
    end
    assign _2997 = { _3860,
                     _326 };
    assign _2994 = { _3860,
                     _316 };
    assign _2991 = { _3860,
                     _276 };
    assign _2988 = { _3860,
                     _271 };
    assign _2986 = { _3860,
                     _266 };
    assign _2989 = _2986 + _2988;
    assign _2992 = _2989 + _2991;
    assign _2995 = _2992 + _2994;
    assign _2998 = _2995 + _2997;
    assign _3001 = _2998 + _3000;
    assign _3004 = _3001 + _3003;
    assign _3007 = _3004 + _3006;
    assign _3009 = _3007 < _3863;
    assign _3010 = _321 & _3009;
    assign _3775 = ~ _3010;
    assign _3776 = _321 & _3775;
    assign _3777 = _213 ? _3776 : _321;
    assign _3778 = _210 ? _316 : _3777;
    assign _182 = _3778;
    always @(posedge _205) begin
        if (_203)
            _321 <= _220;
        else
            _321 <= _182;
    end
    assign _3019 = { _3860,
                     _321 };
    assign _3016 = { _3860,
                     _271 };
    assign _3014 = { _3860,
                     _266 };
    assign _3017 = _3014 + _3016;
    assign _3020 = _3017 + _3019;
    assign _3023 = _3020 + _3022;
    assign _3026 = _3023 + _3025;
    assign _3028 = _3026 < _3863;
    assign _3029 = _316 & _3028;
    assign _3779 = ~ _3029;
    assign _3780 = _316 & _3779;
    assign _3781 = _213 ? _3780 : _316;
    assign _3782 = _210 ? _311 : _3781;
    assign _183 = _3782;
    always @(posedge _205) begin
        if (_203)
            _316 <= _220;
        else
            _316 <= _183;
    end
    assign _3284 = { _3860,
                     _316 };
    assign _3281 = { _3860,
                     _271 };
    assign _3278 = { _3860,
                     _221 };
    assign _3276 = { _3860,
                     _217 };
    assign _3279 = _3276 + _3278;
    assign _3282 = _3279 + _3281;
    assign _3285 = _3282 + _3284;
    assign _3288 = _3285 + _3287;
    assign _3290 = _3288 < _3863;
    assign _3291 = _266 & _3290;
    assign _3783 = ~ _3291;
    assign _3784 = _266 & _3783;
    assign _3785 = _213 ? _3784 : _266;
    assign _3786 = _210 ? _261 : _3785;
    assign _184 = _3786;
    always @(posedge _205) begin
        if (_203)
            _266 <= _220;
        else
            _266 <= _184;
    end
    assign _3256 = { _3860,
                     _266 };
    assign _3253 = { _3860,
                     _226 };
    assign _3250 = { _3860,
                     _221 };
    assign _3248 = { _3860,
                     _217 };
    assign _3251 = _3248 + _3250;
    assign _3254 = _3251 + _3253;
    assign _3257 = _3254 + _3256;
    assign _3260 = _3257 + _3259;
    assign _3263 = _3260 + _3262;
    assign _3266 = _3263 + _3265;
    assign _3269 = _3266 + _3268;
    assign _3271 = _3269 < _3863;
    assign _3272 = _271 & _3271;
    assign _3787 = ~ _3272;
    assign _3788 = _271 & _3787;
    assign _3789 = _213 ? _3788 : _271;
    assign _3790 = _210 ? _266 : _3789;
    assign _185 = _3790;
    always @(posedge _205) begin
        if (_203)
            _271 <= _220;
        else
            _271 <= _185;
    end
    assign _3228 = { _3860,
                     _271 };
    assign _3225 = { _3860,
                     _231 };
    assign _3222 = { _3860,
                     _226 };
    assign _3220 = { _3860,
                     _221 };
    assign _3223 = _3220 + _3222;
    assign _3226 = _3223 + _3225;
    assign _3229 = _3226 + _3228;
    assign _3232 = _3229 + _3231;
    assign _3235 = _3232 + _3234;
    assign _3238 = _3235 + _3237;
    assign _3241 = _3238 + _3240;
    assign _3243 = _3241 < _3863;
    assign _3244 = _276 & _3243;
    assign _3791 = ~ _3244;
    assign _3792 = _276 & _3791;
    assign _3793 = _213 ? _3792 : _276;
    assign _3794 = _210 ? _271 : _3793;
    assign _186 = _3794;
    always @(posedge _205) begin
        if (_203)
            _276 <= _220;
        else
            _276 <= _186;
    end
    assign _3200 = { _3860,
                     _276 };
    assign _3197 = { _3860,
                     _236 };
    assign _3194 = { _3860,
                     _231 };
    assign _3192 = { _3860,
                     _226 };
    assign _3195 = _3192 + _3194;
    assign _3198 = _3195 + _3197;
    assign _3201 = _3198 + _3200;
    assign _3204 = _3201 + _3203;
    assign _3207 = _3204 + _3206;
    assign _3210 = _3207 + _3209;
    assign _3213 = _3210 + _3212;
    assign _3215 = _3213 < _3863;
    assign _3216 = _281 & _3215;
    assign _3795 = ~ _3216;
    assign _3796 = _281 & _3795;
    assign _3797 = _213 ? _3796 : _281;
    assign _3798 = _210 ? _276 : _3797;
    assign _187 = _3798;
    always @(posedge _205) begin
        if (_203)
            _281 <= _220;
        else
            _281 <= _187;
    end
    assign _3172 = { _3860,
                     _281 };
    assign _3169 = { _3860,
                     _241 };
    assign _3166 = { _3860,
                     _236 };
    assign _3164 = { _3860,
                     _231 };
    assign _3167 = _3164 + _3166;
    assign _3170 = _3167 + _3169;
    assign _3173 = _3170 + _3172;
    assign _3176 = _3173 + _3175;
    assign _3179 = _3176 + _3178;
    assign _3182 = _3179 + _3181;
    assign _3185 = _3182 + _3184;
    assign _3187 = _3185 < _3863;
    assign _3188 = _286 & _3187;
    assign _3799 = ~ _3188;
    assign _3800 = _286 & _3799;
    assign _3801 = _213 ? _3800 : _286;
    assign _3802 = _210 ? _281 : _3801;
    assign _188 = _3802;
    always @(posedge _205) begin
        if (_203)
            _286 <= _220;
        else
            _286 <= _188;
    end
    assign _3144 = { _3860,
                     _286 };
    assign _3141 = { _3860,
                     _246 };
    assign _3138 = { _3860,
                     _241 };
    assign _3136 = { _3860,
                     _236 };
    assign _3139 = _3136 + _3138;
    assign _3142 = _3139 + _3141;
    assign _3145 = _3142 + _3144;
    assign _3148 = _3145 + _3147;
    assign _3151 = _3148 + _3150;
    assign _3154 = _3151 + _3153;
    assign _3157 = _3154 + _3156;
    assign _3159 = _3157 < _3863;
    assign _3160 = _291 & _3159;
    assign _3803 = ~ _3160;
    assign _3804 = _291 & _3803;
    assign _3805 = _213 ? _3804 : _291;
    assign _3806 = _210 ? _286 : _3805;
    assign _189 = _3806;
    always @(posedge _205) begin
        if (_203)
            _291 <= _220;
        else
            _291 <= _189;
    end
    assign _3116 = { _3860,
                     _291 };
    assign _3113 = { _3860,
                     _251 };
    assign _3110 = { _3860,
                     _246 };
    assign _3108 = { _3860,
                     _241 };
    assign _3111 = _3108 + _3110;
    assign _3114 = _3111 + _3113;
    assign _3117 = _3114 + _3116;
    assign _3120 = _3117 + _3119;
    assign _3123 = _3120 + _3122;
    assign _3126 = _3123 + _3125;
    assign _3129 = _3126 + _3128;
    assign _3131 = _3129 < _3863;
    assign _3132 = _296 & _3131;
    assign _3807 = ~ _3132;
    assign _3808 = _296 & _3807;
    assign _3809 = _213 ? _3808 : _296;
    assign _3810 = _210 ? _291 : _3809;
    assign _190 = _3810;
    always @(posedge _205) begin
        if (_203)
            _296 <= _220;
        else
            _296 <= _190;
    end
    assign _3088 = { _3860,
                     _296 };
    assign _3085 = { _3860,
                     _256 };
    assign _3082 = { _3860,
                     _251 };
    assign _3080 = { _3860,
                     _246 };
    assign _3083 = _3080 + _3082;
    assign _3086 = _3083 + _3085;
    assign _3089 = _3086 + _3088;
    assign _3092 = _3089 + _3091;
    assign _3095 = _3092 + _3094;
    assign _3098 = _3095 + _3097;
    assign _3101 = _3098 + _3100;
    assign _3103 = _3101 < _3863;
    assign _3104 = _301 & _3103;
    assign _3811 = ~ _3104;
    assign _3812 = _301 & _3811;
    assign _3813 = _213 ? _3812 : _301;
    assign _3814 = _210 ? _296 : _3813;
    assign _191 = _3814;
    always @(posedge _205) begin
        if (_203)
            _301 <= _220;
        else
            _301 <= _191;
    end
    assign _3060 = { _3860,
                     _301 };
    assign _3057 = { _3860,
                     _261 };
    assign _3054 = { _3860,
                     _256 };
    assign _3052 = { _3860,
                     _251 };
    assign _3055 = _3052 + _3054;
    assign _3058 = _3055 + _3057;
    assign _3061 = _3058 + _3060;
    assign _3064 = _3061 + _3063;
    assign _3067 = _3064 + _3066;
    assign _3070 = _3067 + _3069;
    assign _3073 = _3070 + _3072;
    assign _3075 = _3073 < _3863;
    assign _3076 = _306 & _3075;
    assign _3815 = ~ _3076;
    assign _3816 = _306 & _3815;
    assign _3817 = _213 ? _3816 : _306;
    assign _3818 = _210 ? _301 : _3817;
    assign _192 = _3818;
    always @(posedge _205) begin
        if (_203)
            _306 <= _220;
        else
            _306 <= _192;
    end
    assign _3297 = { _3860,
                     _306 };
    assign _3295 = { _3860,
                     _256 };
    assign _3298 = _3295 + _3297;
    assign _3301 = _3298 + _3300;
    assign _3303 = _3301 < _3863;
    assign _3304 = _261 & _3303;
    assign _3819 = ~ _3304;
    assign _3820 = _261 & _3819;
    assign _3821 = _213 ? _3820 : _261;
    assign _3822 = _210 ? _256 : _3821;
    assign _193 = _3822;
    always @(posedge _205) begin
        if (_203)
            _261 <= _220;
        else
            _261 <= _193;
    end
    assign _3310 = { _3860,
                     _261 };
    assign _3308 = { _3860,
                     _251 };
    assign _3311 = _3308 + _3310;
    assign _3314 = _3311 + _3313;
    assign _3317 = _3314 + _3316;
    assign _3320 = _3317 + _3319;
    assign _3322 = _3320 < _3863;
    assign _3323 = _256 & _3322;
    assign _3823 = ~ _3323;
    assign _3824 = _256 & _3823;
    assign _3825 = _213 ? _3824 : _256;
    assign _3826 = _210 ? _251 : _3825;
    assign _194 = _3826;
    always @(posedge _205) begin
        if (_203)
            _256 <= _220;
        else
            _256 <= _194;
    end
    assign _3329 = { _3860,
                     _256 };
    assign _3327 = { _3860,
                     _246 };
    assign _3330 = _3327 + _3329;
    assign _3333 = _3330 + _3332;
    assign _3336 = _3333 + _3335;
    assign _3339 = _3336 + _3338;
    assign _3341 = _3339 < _3863;
    assign _3342 = _251 & _3341;
    assign _3827 = ~ _3342;
    assign _3828 = _251 & _3827;
    assign _3829 = _213 ? _3828 : _251;
    assign _3830 = _210 ? _246 : _3829;
    assign _195 = _3830;
    always @(posedge _205) begin
        if (_203)
            _251 <= _220;
        else
            _251 <= _195;
    end
    assign _3348 = { _3860,
                     _251 };
    assign _3346 = { _3860,
                     _241 };
    assign _3349 = _3346 + _3348;
    assign _3352 = _3349 + _3351;
    assign _3355 = _3352 + _3354;
    assign _3358 = _3355 + _3357;
    assign _3360 = _3358 < _3863;
    assign _3361 = _246 & _3360;
    assign _3831 = ~ _3361;
    assign _3832 = _246 & _3831;
    assign _3833 = _213 ? _3832 : _246;
    assign _3834 = _210 ? _241 : _3833;
    assign _196 = _3834;
    always @(posedge _205) begin
        if (_203)
            _246 <= _220;
        else
            _246 <= _196;
    end
    assign _3367 = { _3860,
                     _246 };
    assign _3365 = { _3860,
                     _236 };
    assign _3368 = _3365 + _3367;
    assign _3371 = _3368 + _3370;
    assign _3374 = _3371 + _3373;
    assign _3377 = _3374 + _3376;
    assign _3379 = _3377 < _3863;
    assign _3380 = _241 & _3379;
    assign _3835 = ~ _3380;
    assign _3836 = _241 & _3835;
    assign _3837 = _213 ? _3836 : _241;
    assign _3838 = _210 ? _236 : _3837;
    assign _197 = _3838;
    always @(posedge _205) begin
        if (_203)
            _241 <= _220;
        else
            _241 <= _197;
    end
    assign _3386 = { _3860,
                     _241 };
    assign _3384 = { _3860,
                     _231 };
    assign _3387 = _3384 + _3386;
    assign _3390 = _3387 + _3389;
    assign _3393 = _3390 + _3392;
    assign _3396 = _3393 + _3395;
    assign _3398 = _3396 < _3863;
    assign _3399 = _236 & _3398;
    assign _3839 = ~ _3399;
    assign _3840 = _236 & _3839;
    assign _3841 = _213 ? _3840 : _236;
    assign _3842 = _210 ? _231 : _3841;
    assign _198 = _3842;
    always @(posedge _205) begin
        if (_203)
            _236 <= _220;
        else
            _236 <= _198;
    end
    assign _3405 = { _3860,
                     _236 };
    assign _3403 = { _3860,
                     _226 };
    assign _3406 = _3403 + _3405;
    assign _3409 = _3406 + _3408;
    assign _3412 = _3409 + _3411;
    assign _3415 = _3412 + _3414;
    assign _3417 = _3415 < _3863;
    assign _3418 = _231 & _3417;
    assign _3843 = ~ _3418;
    assign _3844 = _231 & _3843;
    assign _3845 = _213 ? _3844 : _231;
    assign _3846 = _210 ? _226 : _3845;
    assign _199 = _3846;
    always @(posedge _205) begin
        if (_203)
            _231 <= _220;
        else
            _231 <= _199;
    end
    assign _3424 = { _3860,
                     _231 };
    assign _3422 = { _3860,
                     _221 };
    assign _3425 = _3422 + _3424;
    assign _3428 = _3425 + _3427;
    assign _3431 = _3428 + _3430;
    assign _3434 = _3431 + _3433;
    assign _3436 = _3434 < _3863;
    assign _3437 = _226 & _3436;
    assign _3847 = ~ _3437;
    assign _3848 = _226 & _3847;
    assign _3849 = _213 ? _3848 : _226;
    assign _3850 = _210 ? _221 : _3849;
    assign _200 = _3850;
    always @(posedge _205) begin
        if (_203)
            _226 <= _220;
        else
            _226 <= _200;
    end
    assign _3443 = { _3860,
                     _226 };
    assign _3441 = { _3860,
                     _217 };
    assign _3444 = _3441 + _3443;
    assign _3447 = _3444 + _3446;
    assign _3450 = _3447 + _3449;
    assign _3453 = _3450 + _3452;
    assign _3455 = _3453 < _3863;
    assign _3456 = _221 & _3455;
    assign _3851 = ~ _3456;
    assign _3852 = _221 & _3851;
    assign _3853 = _213 ? _3852 : _221;
    assign _3854 = _210 ? _217 : _3853;
    assign _201 = _3854;
    always @(posedge _205) begin
        if (_203)
            _221 <= _220;
        else
            _221 <= _201;
    end
    assign _3856 = { _3860,
                     _221 };
    assign _3859 = _3856 + _3858;
    assign _3862 = _3859 + _3861;
    assign _3864 = _3862 < _3863;
    assign _203 = clear;
    assign _205 = clock;
    assign _207 = load_data;
    assign _3866 = ~ _3865;
    assign _3867 = _217 & _3866;
    assign _3868 = _213 ? _3867 : _217;
    assign _3869 = _210 ? _207 : _3868;
    assign _208 = _3869;
    always @(posedge _205) begin
        if (_203)
            _217 <= _220;
        else
            _217 <= _208;
    end
    assign _3865 = _217 & _3864;
    assign gnd = 1'b0;
    assign _3870 = _213 ? _3865 : gnd;
    assign _210 = load;
    assign _3871 = _210 ? gnd : _3870;
    assign _211 = _3871;
    assign _719 = { _709,
                    _211 };
    assign _722 = _719 + _721;
    assign _725 = _722 + _724;
    assign _728 = _725 + _727;
    assign _731 = _728 + _730;
    assign _734 = _731 + _733;
    assign _737 = _734 + _736;
    assign _740 = _737 + _739;
    assign _743 = _740 + _742;
    assign _746 = _743 + _745;
    assign _749 = _746 + _748;
    assign _752 = _749 + _751;
    assign _755 = _752 + _754;
    assign _758 = _755 + _757;
    assign _761 = _758 + _760;
    assign _764 = _761 + _763;
    assign _767 = _764 + _766;
    assign _770 = _767 + _769;
    assign _773 = _770 + _772;
    assign _776 = _773 + _775;
    assign _779 = _776 + _778;
    assign _782 = _779 + _781;
    assign _785 = _782 + _784;
    assign _788 = _785 + _787;
    assign _791 = _788 + _790;
    assign _794 = _791 + _793;
    assign _797 = _794 + _796;
    assign _800 = _797 + _799;
    assign _803 = _800 + _802;
    assign _806 = _803 + _805;
    assign _809 = _806 + _808;
    assign _812 = _809 + _811;
    assign _815 = _812 + _814;
    assign _818 = _815 + _817;
    assign _821 = _818 + _820;
    assign _824 = _821 + _823;
    assign _827 = _824 + _826;
    assign _830 = _827 + _829;
    assign _833 = _830 + _832;
    assign _836 = _833 + _835;
    assign _839 = _836 + _838;
    assign _842 = _839 + _841;
    assign _845 = _842 + _844;
    assign _848 = _845 + _847;
    assign _851 = _848 + _850;
    assign _854 = _851 + _853;
    assign _857 = _854 + _856;
    assign _860 = _857 + _859;
    assign _863 = _860 + _862;
    assign _866 = _863 + _865;
    assign _869 = _866 + _868;
    assign _872 = _869 + _871;
    assign _875 = _872 + _874;
    assign _878 = _875 + _877;
    assign _881 = _878 + _880;
    assign _884 = _881 + _883;
    assign _887 = _884 + _886;
    assign _890 = _887 + _889;
    assign _893 = _890 + _892;
    assign _896 = _893 + _895;
    assign _899 = _896 + _898;
    assign _902 = _899 + _901;
    assign _905 = _902 + _904;
    assign _908 = _905 + _907;
    assign _911 = _908 + _910;
    assign _914 = _911 + _913;
    assign _917 = _914 + _916;
    assign _920 = _917 + _919;
    assign _923 = _920 + _922;
    assign _926 = _923 + _925;
    assign _929 = _926 + _928;
    assign _932 = _929 + _931;
    assign _935 = _932 + _934;
    assign _938 = _935 + _937;
    assign _941 = _938 + _940;
    assign _944 = _941 + _943;
    assign _947 = _944 + _946;
    assign _950 = _947 + _949;
    assign _953 = _950 + _952;
    assign _956 = _953 + _955;
    assign _959 = _956 + _958;
    assign _962 = _959 + _961;
    assign _965 = _962 + _964;
    assign _968 = _965 + _967;
    assign _971 = _968 + _970;
    assign _974 = _971 + _973;
    assign _977 = _974 + _976;
    assign _980 = _977 + _979;
    assign _983 = _980 + _982;
    assign _986 = _983 + _985;
    assign _989 = _986 + _988;
    assign _992 = _989 + _991;
    assign _995 = _992 + _994;
    assign _998 = _995 + _997;
    assign _1001 = _998 + _1000;
    assign _1004 = _1001 + _1003;
    assign _1007 = _1004 + _1006;
    assign _1010 = _1007 + _1009;
    assign _1013 = _1010 + _1012;
    assign _1016 = _1013 + _1015;
    assign _3873 = _1016 == _714;
    assign _213 = start;
    assign _3874 = _213 & _3873;
    assign finished = _3874;
    assign total_removed = _715;
    assign current_active = _713;

endmodule
module aoc_solver_top (
    start,
    load_data,
    load,
    clear,
    clock,
    finished,
    total_removed,
    current_active
);

    input start;
    input load_data;
    input load;
    input clear;
    input clock;
    output finished;
    output [15:0] total_removed;
    output [15:0] current_active;

    wire [15:0] _15;
    wire [15:0] _16;
    wire _4;
    wire _6;
    wire _8;
    wire _10;
    wire _12;
    wire [32:0] _14;
    wire _17;
    assign _15 = _14[32:17];
    assign _16 = _14[16:1];
    assign _4 = start;
    assign _6 = load_data;
    assign _8 = load;
    assign _10 = clear;
    assign _12 = clock;
    aoc_solver
        aoc_solver
        ( .clock(_12),
          .clear(_10),
          .load(_8),
          .load_data(_6),
          .start(_4),
          .finished(_14[0:0]),
          .total_removed(_14[16:1]),
          .current_active(_14[32:17]) );
    assign _17 = _14[0:0];
    assign finished = _17;
    assign total_removed = _16;
    assign current_active = _15;

endmodule

