module aoc_solver (
    write_enable,
    clear,
    clock,
    write_data,
    write_addr,
    read_data
);

    input write_enable;
    input clear;
    input clock;
    input [31:0] write_data;
    input [3:0] write_addr;
    output [31:0] read_data;

    wire [14:0] _3889;
    wire [15:0] _3890;
    wire [15:0] _3887;
    wire [15:0] _3884;
    wire [15:0] _3881;
    wire [15:0] _3878;
    wire [15:0] _3875;
    wire [15:0] _3872;
    wire [15:0] _3869;
    wire [15:0] _3866;
    wire [15:0] _3863;
    wire [15:0] _3860;
    wire [15:0] _3857;
    wire [15:0] _3854;
    wire [15:0] _3851;
    wire [15:0] _3848;
    wire [15:0] _3845;
    wire [15:0] _3842;
    wire [15:0] _3839;
    wire [15:0] _3836;
    wire [15:0] _3833;
    wire [15:0] _3830;
    wire [15:0] _3827;
    wire [15:0] _3824;
    wire [15:0] _3821;
    wire [15:0] _3818;
    wire [15:0] _3815;
    wire [15:0] _3812;
    wire [15:0] _3809;
    wire [15:0] _3806;
    wire [15:0] _3803;
    wire [15:0] _3800;
    wire [15:0] _3797;
    wire [15:0] _3794;
    wire [15:0] _3791;
    wire [15:0] _3788;
    wire [15:0] _3785;
    wire [15:0] _3782;
    wire [15:0] _3779;
    wire [15:0] _3776;
    wire [15:0] _3773;
    wire [15:0] _3770;
    wire [15:0] _3767;
    wire [15:0] _3764;
    wire [15:0] _3761;
    wire [15:0] _3758;
    wire [15:0] _3755;
    wire [15:0] _3752;
    wire [15:0] _3749;
    wire [15:0] _3746;
    wire [15:0] _3743;
    wire [15:0] _3740;
    wire [15:0] _3737;
    wire [15:0] _3734;
    wire [15:0] _3731;
    wire [15:0] _3728;
    wire [15:0] _3725;
    wire [15:0] _3722;
    wire [15:0] _3719;
    wire [15:0] _3716;
    wire [15:0] _3713;
    wire [15:0] _3710;
    wire [15:0] _3707;
    wire [15:0] _3704;
    wire [15:0] _3701;
    wire [15:0] _3698;
    wire [15:0] _3695;
    wire [15:0] _3692;
    wire [15:0] _3689;
    wire [15:0] _3686;
    wire [15:0] _3683;
    wire [15:0] _3680;
    wire [15:0] _3677;
    wire [15:0] _3674;
    wire [15:0] _3671;
    wire [15:0] _3668;
    wire [15:0] _3665;
    wire [15:0] _3662;
    wire [15:0] _3659;
    wire [15:0] _3656;
    wire [15:0] _3653;
    wire [15:0] _3650;
    wire [15:0] _3647;
    wire [15:0] _3644;
    wire [15:0] _3641;
    wire [15:0] _3638;
    wire [15:0] _3635;
    wire [15:0] _3632;
    wire [15:0] _3629;
    wire [15:0] _3626;
    wire [15:0] _3623;
    wire [15:0] _3620;
    wire [15:0] _3617;
    wire [15:0] _3614;
    wire [15:0] _3611;
    wire [15:0] _3608;
    wire [15:0] _3605;
    wire [15:0] _3602;
    wire [15:0] _3599;
    wire [15:0] _3596;
    wire [15:0] _3594;
    wire [15:0] _3597;
    wire [15:0] _3600;
    wire [15:0] _3603;
    wire [15:0] _3606;
    wire [15:0] _3609;
    wire [15:0] _3612;
    wire [15:0] _3615;
    wire [15:0] _3618;
    wire [15:0] _3621;
    wire [15:0] _3624;
    wire [15:0] _3627;
    wire [15:0] _3630;
    wire [15:0] _3633;
    wire [15:0] _3636;
    wire [15:0] _3639;
    wire [15:0] _3642;
    wire [15:0] _3645;
    wire [15:0] _3648;
    wire [15:0] _3651;
    wire [15:0] _3654;
    wire [15:0] _3657;
    wire [15:0] _3660;
    wire [15:0] _3663;
    wire [15:0] _3666;
    wire [15:0] _3669;
    wire [15:0] _3672;
    wire [15:0] _3675;
    wire [15:0] _3678;
    wire [15:0] _3681;
    wire [15:0] _3684;
    wire [15:0] _3687;
    wire [15:0] _3690;
    wire [15:0] _3693;
    wire [15:0] _3696;
    wire [15:0] _3699;
    wire [15:0] _3702;
    wire [15:0] _3705;
    wire [15:0] _3708;
    wire [15:0] _3711;
    wire [15:0] _3714;
    wire [15:0] _3717;
    wire [15:0] _3720;
    wire [15:0] _3723;
    wire [15:0] _3726;
    wire [15:0] _3729;
    wire [15:0] _3732;
    wire [15:0] _3735;
    wire [15:0] _3738;
    wire [15:0] _3741;
    wire [15:0] _3744;
    wire [15:0] _3747;
    wire [15:0] _3750;
    wire [15:0] _3753;
    wire [15:0] _3756;
    wire [15:0] _3759;
    wire [15:0] _3762;
    wire [15:0] _3765;
    wire [15:0] _3768;
    wire [15:0] _3771;
    wire [15:0] _3774;
    wire [15:0] _3777;
    wire [15:0] _3780;
    wire [15:0] _3783;
    wire [15:0] _3786;
    wire [15:0] _3789;
    wire [15:0] _3792;
    wire [15:0] _3795;
    wire [15:0] _3798;
    wire [15:0] _3801;
    wire [15:0] _3804;
    wire [15:0] _3807;
    wire [15:0] _3810;
    wire [15:0] _3813;
    wire [15:0] _3816;
    wire [15:0] _3819;
    wire [15:0] _3822;
    wire [15:0] _3825;
    wire [15:0] _3828;
    wire [15:0] _3831;
    wire [15:0] _3834;
    wire [15:0] _3837;
    wire [15:0] _3840;
    wire [15:0] _3843;
    wire [15:0] _3846;
    wire [15:0] _3849;
    wire [15:0] _3852;
    wire [15:0] _3855;
    wire [15:0] _3858;
    wire [15:0] _3861;
    wire [15:0] _3864;
    wire [15:0] _3867;
    wire [15:0] _3870;
    wire [15:0] _3873;
    wire [15:0] _3876;
    wire [15:0] _3879;
    wire [15:0] _3882;
    wire [15:0] _3885;
    wire [15:0] _3888;
    wire [15:0] _3891;
    wire [15:0] _3592;
    wire [31:0] _3892;
    wire [15:0] _525;
    wire [15:0] _225;
    wire [15:0] _526;
    wire [15:0] _1;
    reg [15:0] _223;
    wire [31:0] _3591;
    wire _550;
    wire _551;
    wire _2;
    wire [15:0] _523;
    wire _573;
    wire _574;
    wire _3;
    wire [15:0] _520;
    wire _596;
    wire _597;
    wire _4;
    wire [15:0] _517;
    wire _619;
    wire _620;
    wire _5;
    wire [15:0] _514;
    wire _642;
    wire _643;
    wire _6;
    wire [15:0] _511;
    wire _665;
    wire _666;
    wire _7;
    wire [15:0] _508;
    wire _688;
    wire _689;
    wire _8;
    wire [15:0] _505;
    wire _711;
    wire _712;
    wire _9;
    wire [15:0] _502;
    wire _734;
    wire _735;
    wire _10;
    wire [15:0] _499;
    wire _747;
    wire _748;
    wire _11;
    wire [15:0] _496;
    wire _770;
    wire _771;
    wire _12;
    wire [15:0] _493;
    wire _800;
    wire _801;
    wire _13;
    wire [15:0] _490;
    wire _830;
    wire _831;
    wire _14;
    wire [15:0] _487;
    wire _860;
    wire _861;
    wire _15;
    wire [15:0] _484;
    wire _890;
    wire _891;
    wire _16;
    wire [15:0] _481;
    wire _920;
    wire _921;
    wire _17;
    wire [15:0] _478;
    wire _950;
    wire _951;
    wire _18;
    wire [15:0] _475;
    wire _980;
    wire _981;
    wire _19;
    wire [15:0] _472;
    wire _1010;
    wire _1011;
    wire _20;
    wire [15:0] _469;
    wire _1029;
    wire _1030;
    wire _21;
    wire [15:0] _466;
    wire _1052;
    wire _1053;
    wire _22;
    wire [15:0] _463;
    wire _1082;
    wire _1083;
    wire _23;
    wire [15:0] _460;
    wire _1112;
    wire _1113;
    wire _24;
    wire [15:0] _457;
    wire _1142;
    wire _1143;
    wire _25;
    wire [15:0] _454;
    wire _1172;
    wire _1173;
    wire _26;
    wire [15:0] _451;
    wire _1202;
    wire _1203;
    wire _27;
    wire [15:0] _448;
    wire _1232;
    wire _1233;
    wire _28;
    wire [15:0] _445;
    wire _1262;
    wire _1263;
    wire _29;
    wire [15:0] _442;
    wire _1292;
    wire _1293;
    wire _30;
    wire [15:0] _439;
    wire _1311;
    wire _1312;
    wire _31;
    wire [15:0] _436;
    wire _1334;
    wire _1335;
    wire _32;
    wire [15:0] _433;
    wire _1364;
    wire _1365;
    wire _33;
    wire [15:0] _430;
    wire _1394;
    wire _1395;
    wire _34;
    wire [15:0] _427;
    wire _1424;
    wire _1425;
    wire _35;
    wire [15:0] _424;
    wire _1454;
    wire _1455;
    wire _36;
    wire [15:0] _421;
    wire _1484;
    wire _1485;
    wire _37;
    wire [15:0] _418;
    wire _1514;
    wire _1515;
    wire _38;
    wire [15:0] _415;
    wire _1544;
    wire _1545;
    wire _39;
    wire [15:0] _412;
    wire _1574;
    wire _1575;
    wire _40;
    wire [15:0] _409;
    wire _1593;
    wire _1594;
    wire _41;
    wire [15:0] _406;
    wire _1616;
    wire _1617;
    wire _42;
    wire [15:0] _403;
    wire _1646;
    wire _1647;
    wire _43;
    wire [15:0] _400;
    wire _1676;
    wire _1677;
    wire _44;
    wire [15:0] _397;
    wire _1706;
    wire _1707;
    wire _45;
    wire [15:0] _394;
    wire _1736;
    wire _1737;
    wire _46;
    wire [15:0] _391;
    wire _1766;
    wire _1767;
    wire _47;
    wire [15:0] _388;
    wire _1796;
    wire _1797;
    wire _48;
    wire [15:0] _385;
    wire _1826;
    wire _1827;
    wire _49;
    wire [15:0] _382;
    wire _1856;
    wire _1857;
    wire _50;
    wire [15:0] _379;
    wire _1875;
    wire _1876;
    wire _51;
    wire [15:0] _376;
    wire _1898;
    wire _1899;
    wire _52;
    wire [15:0] _373;
    wire _1928;
    wire _1929;
    wire _53;
    wire [15:0] _370;
    wire _1958;
    wire _1959;
    wire _54;
    wire [15:0] _367;
    wire _1988;
    wire _1989;
    wire _55;
    wire [15:0] _364;
    wire _2018;
    wire _2019;
    wire _56;
    wire [15:0] _361;
    wire _2048;
    wire _2049;
    wire _57;
    wire [15:0] _358;
    wire _2078;
    wire _2079;
    wire _58;
    wire [15:0] _355;
    wire _2108;
    wire _2109;
    wire _59;
    wire [15:0] _352;
    wire _2138;
    wire _2139;
    wire _60;
    wire [15:0] _349;
    wire _2157;
    wire _2158;
    wire _61;
    wire [15:0] _346;
    wire _2180;
    wire _2181;
    wire _62;
    wire [15:0] _343;
    wire _2210;
    wire _2211;
    wire _63;
    wire [15:0] _340;
    wire _2240;
    wire _2241;
    wire _64;
    wire [15:0] _337;
    wire _2270;
    wire _2271;
    wire _65;
    wire [15:0] _334;
    wire _2300;
    wire _2301;
    wire _66;
    wire [15:0] _331;
    wire _2330;
    wire _2331;
    wire _67;
    wire [15:0] _328;
    wire _2360;
    wire _2361;
    wire _68;
    wire [15:0] _325;
    wire _2390;
    wire _2391;
    wire _69;
    wire [15:0] _322;
    wire _2420;
    wire _2421;
    wire _70;
    wire [15:0] _319;
    wire _2439;
    wire _2440;
    wire _71;
    wire [15:0] _316;
    wire _2462;
    wire _2463;
    wire _72;
    wire [15:0] _313;
    wire _2492;
    wire _2493;
    wire _73;
    wire [15:0] _310;
    wire _2522;
    wire _2523;
    wire _74;
    wire [15:0] _307;
    wire _2552;
    wire _2553;
    wire _75;
    wire [15:0] _304;
    wire _2582;
    wire _2583;
    wire _76;
    wire [15:0] _301;
    wire _2612;
    wire _2613;
    wire _77;
    wire [15:0] _298;
    wire _2642;
    wire _2643;
    wire _78;
    wire [15:0] _295;
    wire _2672;
    wire _2673;
    wire _79;
    wire [15:0] _292;
    wire _2702;
    wire _2703;
    wire _80;
    wire [15:0] _289;
    wire _2721;
    wire _2722;
    wire _81;
    wire [15:0] _286;
    wire _2744;
    wire _2745;
    wire _82;
    wire [15:0] _283;
    wire _2774;
    wire _2775;
    wire _83;
    wire [15:0] _280;
    wire _2804;
    wire _2805;
    wire _84;
    wire [15:0] _277;
    wire _2834;
    wire _2835;
    wire _85;
    wire [15:0] _274;
    wire _2864;
    wire _2865;
    wire _86;
    wire [15:0] _271;
    wire _2894;
    wire _2895;
    wire _87;
    wire [15:0] _268;
    wire _2924;
    wire _2925;
    wire _88;
    wire [15:0] _265;
    wire _2954;
    wire _2955;
    wire _89;
    wire [15:0] _262;
    wire _2984;
    wire _2985;
    wire _90;
    wire [15:0] _259;
    wire _3003;
    wire _3004;
    wire _91;
    wire [15:0] _256;
    wire _3016;
    wire _3017;
    wire _92;
    wire [15:0] _253;
    wire _3035;
    wire _3036;
    wire _93;
    wire [15:0] _250;
    wire _3054;
    wire _3055;
    wire _94;
    wire [15:0] _247;
    wire _3073;
    wire _3074;
    wire _95;
    wire [15:0] _244;
    wire _3092;
    wire _3093;
    wire _96;
    wire [15:0] _241;
    wire _3111;
    wire _3112;
    wire _97;
    wire [15:0] _238;
    wire _3130;
    wire _3131;
    wire _98;
    wire [15:0] _235;
    wire _3149;
    wire _3150;
    wire _99;
    wire [15:0] _232;
    wire _3168;
    wire _3169;
    wire _100;
    wire [15:0] _229;
    wire [3:0] _3574;
    wire [2:0] _3571;
    wire [3:0] _3572;
    wire [3:0] _3569;
    wire _2927;
    wire [3:0] _3163;
    wire [3:0] _3160;
    wire [3:0] _3157;
    wire [3:0] _3144;
    wire [3:0] _3141;
    wire [3:0] _3138;
    wire [3:0] _3125;
    wire [3:0] _3122;
    wire [3:0] _3119;
    wire [3:0] _3106;
    wire [3:0] _3103;
    wire [3:0] _3100;
    wire [3:0] _3087;
    wire [3:0] _3084;
    wire [3:0] _3081;
    wire [3:0] _3068;
    wire [3:0] _3065;
    wire [3:0] _3062;
    wire [3:0] _3049;
    wire [3:0] _3046;
    wire [3:0] _3043;
    wire [3:0] _3030;
    wire [3:0] _3027;
    wire [3:0] _3024;
    wire [3:0] _3011;
    wire [3:0] _2769;
    wire [3:0] _2766;
    wire [3:0] _2763;
    wire [3:0] _2760;
    wire [3:0] _2799;
    wire [3:0] _2796;
    wire [3:0] _2793;
    wire [3:0] _2790;
    wire [3:0] _2829;
    wire [3:0] _2826;
    wire [3:0] _2823;
    wire [3:0] _2820;
    wire [3:0] _2859;
    wire [3:0] _2856;
    wire [3:0] _2853;
    wire [3:0] _2850;
    wire [3:0] _2889;
    wire [3:0] _2886;
    wire [3:0] _2883;
    wire [3:0] _2880;
    wire [3:0] _2919;
    wire [3:0] _2916;
    wire [3:0] _2913;
    wire [3:0] _2910;
    wire [3:0] _2949;
    wire [3:0] _2946;
    wire [3:0] _2943;
    wire [3:0] _2940;
    wire [3:0] _2979;
    wire [3:0] _2976;
    wire [3:0] _2973;
    wire [3:0] _2970;
    wire [3:0] _2998;
    wire [3:0] _2716;
    wire [3:0] _2713;
    wire [3:0] _2697;
    wire [3:0] _2694;
    wire [3:0] _2691;
    wire [3:0] _2667;
    wire [3:0] _2664;
    wire [3:0] _2661;
    wire [3:0] _2637;
    wire [3:0] _2634;
    wire [3:0] _2631;
    wire [3:0] _2607;
    wire [3:0] _2604;
    wire [3:0] _2601;
    wire [3:0] _2577;
    wire [3:0] _2574;
    wire [3:0] _2571;
    wire [3:0] _2547;
    wire [3:0] _2544;
    wire [3:0] _2541;
    wire [3:0] _2517;
    wire [3:0] _2514;
    wire [3:0] _2511;
    wire [3:0] _2487;
    wire [3:0] _2484;
    wire [3:0] _2481;
    wire [3:0] _2478;
    wire [3:0] _2475;
    wire [3:0] _2457;
    wire [3:0] _2205;
    wire [3:0] _2202;
    wire [3:0] _2199;
    wire [3:0] _2196;
    wire [3:0] _2235;
    wire [3:0] _2232;
    wire [3:0] _2229;
    wire [3:0] _2226;
    wire [3:0] _2265;
    wire [3:0] _2262;
    wire [3:0] _2259;
    wire [3:0] _2256;
    wire [3:0] _2295;
    wire [3:0] _2292;
    wire [3:0] _2289;
    wire [3:0] _2286;
    wire [3:0] _2325;
    wire [3:0] _2322;
    wire [3:0] _2319;
    wire [3:0] _2316;
    wire [3:0] _2355;
    wire [3:0] _2352;
    wire [3:0] _2349;
    wire [3:0] _2346;
    wire [3:0] _2385;
    wire [3:0] _2382;
    wire [3:0] _2379;
    wire [3:0] _2376;
    wire [3:0] _2415;
    wire [3:0] _2412;
    wire [3:0] _2409;
    wire [3:0] _2406;
    wire [3:0] _2434;
    wire [3:0] _2152;
    wire [3:0] _2149;
    wire [3:0] _2133;
    wire [3:0] _2130;
    wire [3:0] _2127;
    wire [3:0] _2103;
    wire [3:0] _2100;
    wire [3:0] _2097;
    wire [3:0] _2073;
    wire [3:0] _2070;
    wire [3:0] _2067;
    wire [3:0] _2043;
    wire [3:0] _2040;
    wire [3:0] _2037;
    wire [3:0] _2013;
    wire [3:0] _2010;
    wire [3:0] _2007;
    wire [3:0] _1983;
    wire [3:0] _1980;
    wire [3:0] _1977;
    wire [3:0] _1953;
    wire [3:0] _1950;
    wire [3:0] _1947;
    wire [3:0] _1923;
    wire [3:0] _1920;
    wire [3:0] _1917;
    wire [3:0] _1914;
    wire [3:0] _1911;
    wire [3:0] _1893;
    wire [3:0] _1641;
    wire [3:0] _1638;
    wire [3:0] _1635;
    wire [3:0] _1632;
    wire [3:0] _1671;
    wire [3:0] _1668;
    wire [3:0] _1665;
    wire [3:0] _1662;
    wire [3:0] _1701;
    wire [3:0] _1698;
    wire [3:0] _1695;
    wire [3:0] _1692;
    wire [3:0] _1731;
    wire [3:0] _1728;
    wire [3:0] _1725;
    wire [3:0] _1722;
    wire [3:0] _1761;
    wire [3:0] _1758;
    wire [3:0] _1755;
    wire [3:0] _1752;
    wire [3:0] _1791;
    wire [3:0] _1788;
    wire [3:0] _1785;
    wire [3:0] _1782;
    wire [3:0] _1821;
    wire [3:0] _1818;
    wire [3:0] _1815;
    wire [3:0] _1812;
    wire [3:0] _1851;
    wire [3:0] _1848;
    wire [3:0] _1845;
    wire [3:0] _1842;
    wire [3:0] _1870;
    wire [3:0] _1588;
    wire [3:0] _1585;
    wire [3:0] _1569;
    wire [3:0] _1566;
    wire [3:0] _1563;
    wire [3:0] _1539;
    wire [3:0] _1536;
    wire [3:0] _1533;
    wire [3:0] _1509;
    wire [3:0] _1506;
    wire [3:0] _1503;
    wire [3:0] _1479;
    wire [3:0] _1476;
    wire [3:0] _1473;
    wire [3:0] _1449;
    wire [3:0] _1446;
    wire [3:0] _1443;
    wire [3:0] _1419;
    wire [3:0] _1416;
    wire [3:0] _1413;
    wire [3:0] _1389;
    wire [3:0] _1386;
    wire [3:0] _1383;
    wire [3:0] _1359;
    wire [3:0] _1356;
    wire [3:0] _1353;
    wire [3:0] _1350;
    wire [3:0] _1347;
    wire [3:0] _1329;
    wire [3:0] _1077;
    wire [3:0] _1074;
    wire [3:0] _1071;
    wire [3:0] _1068;
    wire [3:0] _1107;
    wire [3:0] _1104;
    wire [3:0] _1101;
    wire [3:0] _1098;
    wire [3:0] _1137;
    wire [3:0] _1134;
    wire [3:0] _1131;
    wire [3:0] _1128;
    wire [3:0] _1167;
    wire [3:0] _1164;
    wire [3:0] _1161;
    wire [3:0] _1158;
    wire [3:0] _1197;
    wire [3:0] _1194;
    wire [3:0] _1191;
    wire [3:0] _1188;
    wire [3:0] _1227;
    wire [3:0] _1224;
    wire [3:0] _1221;
    wire [3:0] _1218;
    wire [3:0] _1257;
    wire [3:0] _1254;
    wire [3:0] _1251;
    wire [3:0] _1248;
    wire [3:0] _1287;
    wire [3:0] _1284;
    wire [3:0] _1281;
    wire [3:0] _1278;
    wire [3:0] _1306;
    wire [3:0] _1024;
    wire [3:0] _1021;
    wire [3:0] _1005;
    wire [3:0] _1002;
    wire [3:0] _999;
    wire [3:0] _975;
    wire [3:0] _972;
    wire [3:0] _969;
    wire [3:0] _945;
    wire [3:0] _942;
    wire [3:0] _939;
    wire [3:0] _915;
    wire [3:0] _912;
    wire [3:0] _909;
    wire [3:0] _885;
    wire [3:0] _882;
    wire [3:0] _879;
    wire [3:0] _855;
    wire [3:0] _852;
    wire [3:0] _849;
    wire [3:0] _825;
    wire [3:0] _822;
    wire [3:0] _819;
    wire [3:0] _795;
    wire [3:0] _792;
    wire [3:0] _789;
    wire [3:0] _786;
    wire [3:0] _783;
    wire [3:0] _765;
    wire [3:0] _545;
    wire [3:0] _540;
    wire [3:0] _536;
    wire [3:0] _541;
    wire [3:0] _546;
    wire _548;
    wire _549;
    wire _3170;
    wire _3171;
    wire _3172;
    wire _3173;
    wire _101;
    reg _532;
    wire [3:0] _568;
    wire [3:0] _591;
    wire [3:0] _614;
    wire [3:0] _637;
    wire [3:0] _660;
    wire [3:0] _683;
    wire [3:0] _706;
    wire [3:0] _729;
    wire [3:0] _742;
    wire [3:0] _739;
    wire [3:0] _737;
    wire [3:0] _740;
    wire [3:0] _743;
    wire _745;
    wire _746;
    wire _3174;
    wire _3175;
    wire _3176;
    wire _3177;
    wire _102;
    reg _725;
    wire [3:0] _726;
    wire [3:0] _721;
    wire [3:0] _718;
    wire [3:0] _716;
    wire [3:0] _719;
    wire [3:0] _722;
    wire [3:0] _727;
    wire [3:0] _730;
    wire _732;
    wire _733;
    wire _3178;
    wire _3179;
    wire _3180;
    wire _3181;
    wire _103;
    reg _702;
    wire [3:0] _703;
    wire [3:0] _698;
    wire [3:0] _695;
    wire [3:0] _693;
    wire [3:0] _696;
    wire [3:0] _699;
    wire [3:0] _704;
    wire [3:0] _707;
    wire _709;
    wire _710;
    wire _3182;
    wire _3183;
    wire _3184;
    wire _3185;
    wire _104;
    reg _679;
    wire [3:0] _680;
    wire [3:0] _675;
    wire [3:0] _672;
    wire [3:0] _670;
    wire [3:0] _673;
    wire [3:0] _676;
    wire [3:0] _681;
    wire [3:0] _684;
    wire _686;
    wire _687;
    wire _3186;
    wire _3187;
    wire _3188;
    wire _3189;
    wire _105;
    reg _656;
    wire [3:0] _657;
    wire [3:0] _652;
    wire [3:0] _649;
    wire [3:0] _647;
    wire [3:0] _650;
    wire [3:0] _653;
    wire [3:0] _658;
    wire [3:0] _661;
    wire _663;
    wire _664;
    wire _3190;
    wire _3191;
    wire _3192;
    wire _3193;
    wire _106;
    reg _633;
    wire [3:0] _634;
    wire [3:0] _629;
    wire [3:0] _626;
    wire [3:0] _624;
    wire [3:0] _627;
    wire [3:0] _630;
    wire [3:0] _635;
    wire [3:0] _638;
    wire _640;
    wire _641;
    wire _3194;
    wire _3195;
    wire _3196;
    wire _3197;
    wire _107;
    reg _610;
    wire [3:0] _611;
    wire [3:0] _606;
    wire [3:0] _603;
    wire [3:0] _601;
    wire [3:0] _604;
    wire [3:0] _607;
    wire [3:0] _612;
    wire [3:0] _615;
    wire _617;
    wire _618;
    wire _3198;
    wire _3199;
    wire _3200;
    wire _3201;
    wire _108;
    reg _587;
    wire [3:0] _588;
    wire [3:0] _583;
    wire [3:0] _580;
    wire [3:0] _578;
    wire [3:0] _581;
    wire [3:0] _584;
    wire [3:0] _589;
    wire [3:0] _592;
    wire _594;
    wire _595;
    wire _3202;
    wire _3203;
    wire _3204;
    wire _3205;
    wire _109;
    reg _564;
    wire [3:0] _565;
    wire [3:0] _560;
    wire [3:0] _557;
    wire [3:0] _555;
    wire [3:0] _558;
    wire [3:0] _561;
    wire [3:0] _566;
    wire [3:0] _569;
    wire _571;
    wire _572;
    wire _3206;
    wire _3207;
    wire _3208;
    wire _3209;
    wire _110;
    reg _544;
    wire [3:0] _762;
    wire [3:0] _759;
    wire [3:0] _756;
    wire [3:0] _752;
    wire [3:0] _757;
    wire [3:0] _760;
    wire [3:0] _763;
    wire [3:0] _766;
    wire _768;
    wire _769;
    wire _3210;
    wire _3211;
    wire _3212;
    wire _3213;
    wire _111;
    reg _539;
    wire [3:0] _1047;
    wire [3:0] _1044;
    wire [3:0] _1041;
    wire [3:0] _1038;
    wire [3:0] _1034;
    wire [3:0] _1039;
    wire [3:0] _1042;
    wire [3:0] _1045;
    wire [3:0] _1048;
    wire _1050;
    wire _1051;
    wire _3214;
    wire _3215;
    wire _3216;
    wire _3217;
    wire _112;
    reg _755;
    wire [3:0] _780;
    wire [3:0] _777;
    wire [3:0] _775;
    wire [3:0] _778;
    wire [3:0] _781;
    wire [3:0] _784;
    wire [3:0] _787;
    wire [3:0] _790;
    wire [3:0] _793;
    wire [3:0] _796;
    wire _798;
    wire _799;
    wire _3218;
    wire _3219;
    wire _3220;
    wire _3221;
    wire _113;
    reg _535;
    wire [3:0] _816;
    wire [3:0] _813;
    wire [3:0] _810;
    wire [3:0] _807;
    wire [3:0] _805;
    wire [3:0] _808;
    wire [3:0] _811;
    wire [3:0] _814;
    wire [3:0] _817;
    wire [3:0] _820;
    wire [3:0] _823;
    wire [3:0] _826;
    wire _828;
    wire _829;
    wire _3222;
    wire _3223;
    wire _3224;
    wire _3225;
    wire _114;
    reg _554;
    wire [3:0] _846;
    wire [3:0] _843;
    wire [3:0] _840;
    wire [3:0] _837;
    wire [3:0] _835;
    wire [3:0] _838;
    wire [3:0] _841;
    wire [3:0] _844;
    wire [3:0] _847;
    wire [3:0] _850;
    wire [3:0] _853;
    wire [3:0] _856;
    wire _858;
    wire _859;
    wire _3226;
    wire _3227;
    wire _3228;
    wire _3229;
    wire _115;
    reg _577;
    wire [3:0] _876;
    wire [3:0] _873;
    wire [3:0] _870;
    wire [3:0] _867;
    wire [3:0] _865;
    wire [3:0] _868;
    wire [3:0] _871;
    wire [3:0] _874;
    wire [3:0] _877;
    wire [3:0] _880;
    wire [3:0] _883;
    wire [3:0] _886;
    wire _888;
    wire _889;
    wire _3230;
    wire _3231;
    wire _3232;
    wire _3233;
    wire _116;
    reg _600;
    wire [3:0] _906;
    wire [3:0] _903;
    wire [3:0] _900;
    wire [3:0] _897;
    wire [3:0] _895;
    wire [3:0] _898;
    wire [3:0] _901;
    wire [3:0] _904;
    wire [3:0] _907;
    wire [3:0] _910;
    wire [3:0] _913;
    wire [3:0] _916;
    wire _918;
    wire _919;
    wire _3234;
    wire _3235;
    wire _3236;
    wire _3237;
    wire _117;
    reg _623;
    wire [3:0] _936;
    wire [3:0] _933;
    wire [3:0] _930;
    wire [3:0] _927;
    wire [3:0] _925;
    wire [3:0] _928;
    wire [3:0] _931;
    wire [3:0] _934;
    wire [3:0] _937;
    wire [3:0] _940;
    wire [3:0] _943;
    wire [3:0] _946;
    wire _948;
    wire _949;
    wire _3238;
    wire _3239;
    wire _3240;
    wire _3241;
    wire _118;
    reg _646;
    wire [3:0] _966;
    wire [3:0] _963;
    wire [3:0] _960;
    wire [3:0] _957;
    wire [3:0] _955;
    wire [3:0] _958;
    wire [3:0] _961;
    wire [3:0] _964;
    wire [3:0] _967;
    wire [3:0] _970;
    wire [3:0] _973;
    wire [3:0] _976;
    wire _978;
    wire _979;
    wire _3242;
    wire _3243;
    wire _3244;
    wire _3245;
    wire _119;
    reg _669;
    wire [3:0] _996;
    wire [3:0] _993;
    wire [3:0] _990;
    wire [3:0] _987;
    wire [3:0] _985;
    wire [3:0] _988;
    wire [3:0] _991;
    wire [3:0] _994;
    wire [3:0] _997;
    wire [3:0] _1000;
    wire [3:0] _1003;
    wire [3:0] _1006;
    wire _1008;
    wire _1009;
    wire _3246;
    wire _3247;
    wire _3248;
    wire _3249;
    wire _120;
    reg _692;
    wire [3:0] _1018;
    wire [3:0] _1015;
    wire [3:0] _1013;
    wire [3:0] _1016;
    wire [3:0] _1019;
    wire [3:0] _1022;
    wire [3:0] _1025;
    wire _1027;
    wire _1028;
    wire _3250;
    wire _3251;
    wire _3252;
    wire _3253;
    wire _121;
    reg _715;
    wire [3:0] _1303;
    wire [3:0] _1300;
    wire [3:0] _1297;
    wire [3:0] _1295;
    wire [3:0] _1298;
    wire [3:0] _1301;
    wire [3:0] _1304;
    wire [3:0] _1307;
    wire _1309;
    wire _1310;
    wire _3254;
    wire _3255;
    wire _3256;
    wire _3257;
    wire _122;
    reg _984;
    wire [3:0] _1275;
    wire [3:0] _1272;
    wire [3:0] _1269;
    wire [3:0] _1267;
    wire [3:0] _1270;
    wire [3:0] _1273;
    wire [3:0] _1276;
    wire [3:0] _1279;
    wire [3:0] _1282;
    wire [3:0] _1285;
    wire [3:0] _1288;
    wire _1290;
    wire _1291;
    wire _3258;
    wire _3259;
    wire _3260;
    wire _3261;
    wire _123;
    reg _954;
    wire [3:0] _1245;
    wire [3:0] _1242;
    wire [3:0] _1239;
    wire [3:0] _1237;
    wire [3:0] _1240;
    wire [3:0] _1243;
    wire [3:0] _1246;
    wire [3:0] _1249;
    wire [3:0] _1252;
    wire [3:0] _1255;
    wire [3:0] _1258;
    wire _1260;
    wire _1261;
    wire _3262;
    wire _3263;
    wire _3264;
    wire _3265;
    wire _124;
    reg _924;
    wire [3:0] _1215;
    wire [3:0] _1212;
    wire [3:0] _1209;
    wire [3:0] _1207;
    wire [3:0] _1210;
    wire [3:0] _1213;
    wire [3:0] _1216;
    wire [3:0] _1219;
    wire [3:0] _1222;
    wire [3:0] _1225;
    wire [3:0] _1228;
    wire _1230;
    wire _1231;
    wire _3266;
    wire _3267;
    wire _3268;
    wire _3269;
    wire _125;
    reg _894;
    wire [3:0] _1185;
    wire [3:0] _1182;
    wire [3:0] _1179;
    wire [3:0] _1177;
    wire [3:0] _1180;
    wire [3:0] _1183;
    wire [3:0] _1186;
    wire [3:0] _1189;
    wire [3:0] _1192;
    wire [3:0] _1195;
    wire [3:0] _1198;
    wire _1200;
    wire _1201;
    wire _3270;
    wire _3271;
    wire _3272;
    wire _3273;
    wire _126;
    reg _864;
    wire [3:0] _1155;
    wire [3:0] _1152;
    wire [3:0] _1149;
    wire [3:0] _1147;
    wire [3:0] _1150;
    wire [3:0] _1153;
    wire [3:0] _1156;
    wire [3:0] _1159;
    wire [3:0] _1162;
    wire [3:0] _1165;
    wire [3:0] _1168;
    wire _1170;
    wire _1171;
    wire _3274;
    wire _3275;
    wire _3276;
    wire _3277;
    wire _127;
    reg _834;
    wire [3:0] _1125;
    wire [3:0] _1122;
    wire [3:0] _1119;
    wire [3:0] _1117;
    wire [3:0] _1120;
    wire [3:0] _1123;
    wire [3:0] _1126;
    wire [3:0] _1129;
    wire [3:0] _1132;
    wire [3:0] _1135;
    wire [3:0] _1138;
    wire _1140;
    wire _1141;
    wire _3278;
    wire _3279;
    wire _3280;
    wire _3281;
    wire _128;
    reg _804;
    wire [3:0] _1095;
    wire [3:0] _1092;
    wire [3:0] _1089;
    wire [3:0] _1087;
    wire [3:0] _1090;
    wire [3:0] _1093;
    wire [3:0] _1096;
    wire [3:0] _1099;
    wire [3:0] _1102;
    wire [3:0] _1105;
    wire [3:0] _1108;
    wire _1110;
    wire _1111;
    wire _3282;
    wire _3283;
    wire _3284;
    wire _3285;
    wire _129;
    reg _774;
    wire [3:0] _1065;
    wire [3:0] _1062;
    wire [3:0] _1059;
    wire [3:0] _1057;
    wire [3:0] _1060;
    wire [3:0] _1063;
    wire [3:0] _1066;
    wire [3:0] _1069;
    wire [3:0] _1072;
    wire [3:0] _1075;
    wire [3:0] _1078;
    wire _1080;
    wire _1081;
    wire _3286;
    wire _3287;
    wire _3288;
    wire _3289;
    wire _130;
    reg _751;
    wire [3:0] _1326;
    wire [3:0] _1323;
    wire [3:0] _1320;
    wire [3:0] _1316;
    wire [3:0] _1321;
    wire [3:0] _1324;
    wire [3:0] _1327;
    wire [3:0] _1330;
    wire _1332;
    wire _1333;
    wire _3290;
    wire _3291;
    wire _3292;
    wire _3293;
    wire _131;
    reg _1037;
    wire [3:0] _1611;
    wire [3:0] _1608;
    wire [3:0] _1605;
    wire [3:0] _1602;
    wire [3:0] _1598;
    wire [3:0] _1603;
    wire [3:0] _1606;
    wire [3:0] _1609;
    wire [3:0] _1612;
    wire _1614;
    wire _1615;
    wire _3294;
    wire _3295;
    wire _3296;
    wire _3297;
    wire _132;
    reg _1319;
    wire [3:0] _1344;
    wire [3:0] _1341;
    wire [3:0] _1339;
    wire [3:0] _1342;
    wire [3:0] _1345;
    wire [3:0] _1348;
    wire [3:0] _1351;
    wire [3:0] _1354;
    wire [3:0] _1357;
    wire [3:0] _1360;
    wire _1362;
    wire _1363;
    wire _3298;
    wire _3299;
    wire _3300;
    wire _3301;
    wire _133;
    reg _1033;
    wire [3:0] _1380;
    wire [3:0] _1377;
    wire [3:0] _1374;
    wire [3:0] _1371;
    wire [3:0] _1369;
    wire [3:0] _1372;
    wire [3:0] _1375;
    wire [3:0] _1378;
    wire [3:0] _1381;
    wire [3:0] _1384;
    wire [3:0] _1387;
    wire [3:0] _1390;
    wire _1392;
    wire _1393;
    wire _3302;
    wire _3303;
    wire _3304;
    wire _3305;
    wire _134;
    reg _1056;
    wire [3:0] _1410;
    wire [3:0] _1407;
    wire [3:0] _1404;
    wire [3:0] _1401;
    wire [3:0] _1399;
    wire [3:0] _1402;
    wire [3:0] _1405;
    wire [3:0] _1408;
    wire [3:0] _1411;
    wire [3:0] _1414;
    wire [3:0] _1417;
    wire [3:0] _1420;
    wire _1422;
    wire _1423;
    wire _3306;
    wire _3307;
    wire _3308;
    wire _3309;
    wire _135;
    reg _1086;
    wire [3:0] _1440;
    wire [3:0] _1437;
    wire [3:0] _1434;
    wire [3:0] _1431;
    wire [3:0] _1429;
    wire [3:0] _1432;
    wire [3:0] _1435;
    wire [3:0] _1438;
    wire [3:0] _1441;
    wire [3:0] _1444;
    wire [3:0] _1447;
    wire [3:0] _1450;
    wire _1452;
    wire _1453;
    wire _3310;
    wire _3311;
    wire _3312;
    wire _3313;
    wire _136;
    reg _1116;
    wire [3:0] _1470;
    wire [3:0] _1467;
    wire [3:0] _1464;
    wire [3:0] _1461;
    wire [3:0] _1459;
    wire [3:0] _1462;
    wire [3:0] _1465;
    wire [3:0] _1468;
    wire [3:0] _1471;
    wire [3:0] _1474;
    wire [3:0] _1477;
    wire [3:0] _1480;
    wire _1482;
    wire _1483;
    wire _3314;
    wire _3315;
    wire _3316;
    wire _3317;
    wire _137;
    reg _1146;
    wire [3:0] _1500;
    wire [3:0] _1497;
    wire [3:0] _1494;
    wire [3:0] _1491;
    wire [3:0] _1489;
    wire [3:0] _1492;
    wire [3:0] _1495;
    wire [3:0] _1498;
    wire [3:0] _1501;
    wire [3:0] _1504;
    wire [3:0] _1507;
    wire [3:0] _1510;
    wire _1512;
    wire _1513;
    wire _3318;
    wire _3319;
    wire _3320;
    wire _3321;
    wire _138;
    reg _1176;
    wire [3:0] _1530;
    wire [3:0] _1527;
    wire [3:0] _1524;
    wire [3:0] _1521;
    wire [3:0] _1519;
    wire [3:0] _1522;
    wire [3:0] _1525;
    wire [3:0] _1528;
    wire [3:0] _1531;
    wire [3:0] _1534;
    wire [3:0] _1537;
    wire [3:0] _1540;
    wire _1542;
    wire _1543;
    wire _3322;
    wire _3323;
    wire _3324;
    wire _3325;
    wire _139;
    reg _1206;
    wire [3:0] _1560;
    wire [3:0] _1557;
    wire [3:0] _1554;
    wire [3:0] _1551;
    wire [3:0] _1549;
    wire [3:0] _1552;
    wire [3:0] _1555;
    wire [3:0] _1558;
    wire [3:0] _1561;
    wire [3:0] _1564;
    wire [3:0] _1567;
    wire [3:0] _1570;
    wire _1572;
    wire _1573;
    wire _3326;
    wire _3327;
    wire _3328;
    wire _3329;
    wire _140;
    reg _1236;
    wire [3:0] _1582;
    wire [3:0] _1579;
    wire [3:0] _1577;
    wire [3:0] _1580;
    wire [3:0] _1583;
    wire [3:0] _1586;
    wire [3:0] _1589;
    wire _1591;
    wire _1592;
    wire _3330;
    wire _3331;
    wire _3332;
    wire _3333;
    wire _141;
    reg _1266;
    wire [3:0] _1867;
    wire [3:0] _1864;
    wire [3:0] _1861;
    wire [3:0] _1859;
    wire [3:0] _1862;
    wire [3:0] _1865;
    wire [3:0] _1868;
    wire [3:0] _1871;
    wire _1873;
    wire _1874;
    wire _3334;
    wire _3335;
    wire _3336;
    wire _3337;
    wire _142;
    reg _1548;
    wire [3:0] _1839;
    wire [3:0] _1836;
    wire [3:0] _1833;
    wire [3:0] _1831;
    wire [3:0] _1834;
    wire [3:0] _1837;
    wire [3:0] _1840;
    wire [3:0] _1843;
    wire [3:0] _1846;
    wire [3:0] _1849;
    wire [3:0] _1852;
    wire _1854;
    wire _1855;
    wire _3338;
    wire _3339;
    wire _3340;
    wire _3341;
    wire _143;
    reg _1518;
    wire [3:0] _1809;
    wire [3:0] _1806;
    wire [3:0] _1803;
    wire [3:0] _1801;
    wire [3:0] _1804;
    wire [3:0] _1807;
    wire [3:0] _1810;
    wire [3:0] _1813;
    wire [3:0] _1816;
    wire [3:0] _1819;
    wire [3:0] _1822;
    wire _1824;
    wire _1825;
    wire _3342;
    wire _3343;
    wire _3344;
    wire _3345;
    wire _144;
    reg _1488;
    wire [3:0] _1779;
    wire [3:0] _1776;
    wire [3:0] _1773;
    wire [3:0] _1771;
    wire [3:0] _1774;
    wire [3:0] _1777;
    wire [3:0] _1780;
    wire [3:0] _1783;
    wire [3:0] _1786;
    wire [3:0] _1789;
    wire [3:0] _1792;
    wire _1794;
    wire _1795;
    wire _3346;
    wire _3347;
    wire _3348;
    wire _3349;
    wire _145;
    reg _1458;
    wire [3:0] _1749;
    wire [3:0] _1746;
    wire [3:0] _1743;
    wire [3:0] _1741;
    wire [3:0] _1744;
    wire [3:0] _1747;
    wire [3:0] _1750;
    wire [3:0] _1753;
    wire [3:0] _1756;
    wire [3:0] _1759;
    wire [3:0] _1762;
    wire _1764;
    wire _1765;
    wire _3350;
    wire _3351;
    wire _3352;
    wire _3353;
    wire _146;
    reg _1428;
    wire [3:0] _1719;
    wire [3:0] _1716;
    wire [3:0] _1713;
    wire [3:0] _1711;
    wire [3:0] _1714;
    wire [3:0] _1717;
    wire [3:0] _1720;
    wire [3:0] _1723;
    wire [3:0] _1726;
    wire [3:0] _1729;
    wire [3:0] _1732;
    wire _1734;
    wire _1735;
    wire _3354;
    wire _3355;
    wire _3356;
    wire _3357;
    wire _147;
    reg _1398;
    wire [3:0] _1689;
    wire [3:0] _1686;
    wire [3:0] _1683;
    wire [3:0] _1681;
    wire [3:0] _1684;
    wire [3:0] _1687;
    wire [3:0] _1690;
    wire [3:0] _1693;
    wire [3:0] _1696;
    wire [3:0] _1699;
    wire [3:0] _1702;
    wire _1704;
    wire _1705;
    wire _3358;
    wire _3359;
    wire _3360;
    wire _3361;
    wire _148;
    reg _1368;
    wire [3:0] _1659;
    wire [3:0] _1656;
    wire [3:0] _1653;
    wire [3:0] _1651;
    wire [3:0] _1654;
    wire [3:0] _1657;
    wire [3:0] _1660;
    wire [3:0] _1663;
    wire [3:0] _1666;
    wire [3:0] _1669;
    wire [3:0] _1672;
    wire _1674;
    wire _1675;
    wire _3362;
    wire _3363;
    wire _3364;
    wire _3365;
    wire _149;
    reg _1338;
    wire [3:0] _1629;
    wire [3:0] _1626;
    wire [3:0] _1623;
    wire [3:0] _1621;
    wire [3:0] _1624;
    wire [3:0] _1627;
    wire [3:0] _1630;
    wire [3:0] _1633;
    wire [3:0] _1636;
    wire [3:0] _1639;
    wire [3:0] _1642;
    wire _1644;
    wire _1645;
    wire _3366;
    wire _3367;
    wire _3368;
    wire _3369;
    wire _150;
    reg _1315;
    wire [3:0] _1890;
    wire [3:0] _1887;
    wire [3:0] _1884;
    wire [3:0] _1880;
    wire [3:0] _1885;
    wire [3:0] _1888;
    wire [3:0] _1891;
    wire [3:0] _1894;
    wire _1896;
    wire _1897;
    wire _3370;
    wire _3371;
    wire _3372;
    wire _3373;
    wire _151;
    reg _1601;
    wire [3:0] _2175;
    wire [3:0] _2172;
    wire [3:0] _2169;
    wire [3:0] _2166;
    wire [3:0] _2162;
    wire [3:0] _2167;
    wire [3:0] _2170;
    wire [3:0] _2173;
    wire [3:0] _2176;
    wire _2178;
    wire _2179;
    wire _3374;
    wire _3375;
    wire _3376;
    wire _3377;
    wire _152;
    reg _1883;
    wire [3:0] _1908;
    wire [3:0] _1905;
    wire [3:0] _1903;
    wire [3:0] _1906;
    wire [3:0] _1909;
    wire [3:0] _1912;
    wire [3:0] _1915;
    wire [3:0] _1918;
    wire [3:0] _1921;
    wire [3:0] _1924;
    wire _1926;
    wire _1927;
    wire _3378;
    wire _3379;
    wire _3380;
    wire _3381;
    wire _153;
    reg _1597;
    wire [3:0] _1944;
    wire [3:0] _1941;
    wire [3:0] _1938;
    wire [3:0] _1935;
    wire [3:0] _1933;
    wire [3:0] _1936;
    wire [3:0] _1939;
    wire [3:0] _1942;
    wire [3:0] _1945;
    wire [3:0] _1948;
    wire [3:0] _1951;
    wire [3:0] _1954;
    wire _1956;
    wire _1957;
    wire _3382;
    wire _3383;
    wire _3384;
    wire _3385;
    wire _154;
    reg _1620;
    wire [3:0] _1974;
    wire [3:0] _1971;
    wire [3:0] _1968;
    wire [3:0] _1965;
    wire [3:0] _1963;
    wire [3:0] _1966;
    wire [3:0] _1969;
    wire [3:0] _1972;
    wire [3:0] _1975;
    wire [3:0] _1978;
    wire [3:0] _1981;
    wire [3:0] _1984;
    wire _1986;
    wire _1987;
    wire _3386;
    wire _3387;
    wire _3388;
    wire _3389;
    wire _155;
    reg _1650;
    wire [3:0] _2004;
    wire [3:0] _2001;
    wire [3:0] _1998;
    wire [3:0] _1995;
    wire [3:0] _1993;
    wire [3:0] _1996;
    wire [3:0] _1999;
    wire [3:0] _2002;
    wire [3:0] _2005;
    wire [3:0] _2008;
    wire [3:0] _2011;
    wire [3:0] _2014;
    wire _2016;
    wire _2017;
    wire _3390;
    wire _3391;
    wire _3392;
    wire _3393;
    wire _156;
    reg _1680;
    wire [3:0] _2034;
    wire [3:0] _2031;
    wire [3:0] _2028;
    wire [3:0] _2025;
    wire [3:0] _2023;
    wire [3:0] _2026;
    wire [3:0] _2029;
    wire [3:0] _2032;
    wire [3:0] _2035;
    wire [3:0] _2038;
    wire [3:0] _2041;
    wire [3:0] _2044;
    wire _2046;
    wire _2047;
    wire _3394;
    wire _3395;
    wire _3396;
    wire _3397;
    wire _157;
    reg _1710;
    wire [3:0] _2064;
    wire [3:0] _2061;
    wire [3:0] _2058;
    wire [3:0] _2055;
    wire [3:0] _2053;
    wire [3:0] _2056;
    wire [3:0] _2059;
    wire [3:0] _2062;
    wire [3:0] _2065;
    wire [3:0] _2068;
    wire [3:0] _2071;
    wire [3:0] _2074;
    wire _2076;
    wire _2077;
    wire _3398;
    wire _3399;
    wire _3400;
    wire _3401;
    wire _158;
    reg _1740;
    wire [3:0] _2094;
    wire [3:0] _2091;
    wire [3:0] _2088;
    wire [3:0] _2085;
    wire [3:0] _2083;
    wire [3:0] _2086;
    wire [3:0] _2089;
    wire [3:0] _2092;
    wire [3:0] _2095;
    wire [3:0] _2098;
    wire [3:0] _2101;
    wire [3:0] _2104;
    wire _2106;
    wire _2107;
    wire _3402;
    wire _3403;
    wire _3404;
    wire _3405;
    wire _159;
    reg _1770;
    wire [3:0] _2124;
    wire [3:0] _2121;
    wire [3:0] _2118;
    wire [3:0] _2115;
    wire [3:0] _2113;
    wire [3:0] _2116;
    wire [3:0] _2119;
    wire [3:0] _2122;
    wire [3:0] _2125;
    wire [3:0] _2128;
    wire [3:0] _2131;
    wire [3:0] _2134;
    wire _2136;
    wire _2137;
    wire _3406;
    wire _3407;
    wire _3408;
    wire _3409;
    wire _160;
    reg _1800;
    wire [3:0] _2146;
    wire [3:0] _2143;
    wire [3:0] _2141;
    wire [3:0] _2144;
    wire [3:0] _2147;
    wire [3:0] _2150;
    wire [3:0] _2153;
    wire _2155;
    wire _2156;
    wire _3410;
    wire _3411;
    wire _3412;
    wire _3413;
    wire _161;
    reg _1830;
    wire [3:0] _2431;
    wire [3:0] _2428;
    wire [3:0] _2425;
    wire [3:0] _2423;
    wire [3:0] _2426;
    wire [3:0] _2429;
    wire [3:0] _2432;
    wire [3:0] _2435;
    wire _2437;
    wire _2438;
    wire _3414;
    wire _3415;
    wire _3416;
    wire _3417;
    wire _162;
    reg _2112;
    wire [3:0] _2403;
    wire [3:0] _2400;
    wire [3:0] _2397;
    wire [3:0] _2395;
    wire [3:0] _2398;
    wire [3:0] _2401;
    wire [3:0] _2404;
    wire [3:0] _2407;
    wire [3:0] _2410;
    wire [3:0] _2413;
    wire [3:0] _2416;
    wire _2418;
    wire _2419;
    wire _3418;
    wire _3419;
    wire _3420;
    wire _3421;
    wire _163;
    reg _2082;
    wire [3:0] _2373;
    wire [3:0] _2370;
    wire [3:0] _2367;
    wire [3:0] _2365;
    wire [3:0] _2368;
    wire [3:0] _2371;
    wire [3:0] _2374;
    wire [3:0] _2377;
    wire [3:0] _2380;
    wire [3:0] _2383;
    wire [3:0] _2386;
    wire _2388;
    wire _2389;
    wire _3422;
    wire _3423;
    wire _3424;
    wire _3425;
    wire _164;
    reg _2052;
    wire [3:0] _2343;
    wire [3:0] _2340;
    wire [3:0] _2337;
    wire [3:0] _2335;
    wire [3:0] _2338;
    wire [3:0] _2341;
    wire [3:0] _2344;
    wire [3:0] _2347;
    wire [3:0] _2350;
    wire [3:0] _2353;
    wire [3:0] _2356;
    wire _2358;
    wire _2359;
    wire _3426;
    wire _3427;
    wire _3428;
    wire _3429;
    wire _165;
    reg _2022;
    wire [3:0] _2313;
    wire [3:0] _2310;
    wire [3:0] _2307;
    wire [3:0] _2305;
    wire [3:0] _2308;
    wire [3:0] _2311;
    wire [3:0] _2314;
    wire [3:0] _2317;
    wire [3:0] _2320;
    wire [3:0] _2323;
    wire [3:0] _2326;
    wire _2328;
    wire _2329;
    wire _3430;
    wire _3431;
    wire _3432;
    wire _3433;
    wire _166;
    reg _1992;
    wire [3:0] _2283;
    wire [3:0] _2280;
    wire [3:0] _2277;
    wire [3:0] _2275;
    wire [3:0] _2278;
    wire [3:0] _2281;
    wire [3:0] _2284;
    wire [3:0] _2287;
    wire [3:0] _2290;
    wire [3:0] _2293;
    wire [3:0] _2296;
    wire _2298;
    wire _2299;
    wire _3434;
    wire _3435;
    wire _3436;
    wire _3437;
    wire _167;
    reg _1962;
    wire [3:0] _2253;
    wire [3:0] _2250;
    wire [3:0] _2247;
    wire [3:0] _2245;
    wire [3:0] _2248;
    wire [3:0] _2251;
    wire [3:0] _2254;
    wire [3:0] _2257;
    wire [3:0] _2260;
    wire [3:0] _2263;
    wire [3:0] _2266;
    wire _2268;
    wire _2269;
    wire _3438;
    wire _3439;
    wire _3440;
    wire _3441;
    wire _168;
    reg _1932;
    wire [3:0] _2223;
    wire [3:0] _2220;
    wire [3:0] _2217;
    wire [3:0] _2215;
    wire [3:0] _2218;
    wire [3:0] _2221;
    wire [3:0] _2224;
    wire [3:0] _2227;
    wire [3:0] _2230;
    wire [3:0] _2233;
    wire [3:0] _2236;
    wire _2238;
    wire _2239;
    wire _3442;
    wire _3443;
    wire _3444;
    wire _3445;
    wire _169;
    reg _1902;
    wire [3:0] _2193;
    wire [3:0] _2190;
    wire [3:0] _2187;
    wire [3:0] _2185;
    wire [3:0] _2188;
    wire [3:0] _2191;
    wire [3:0] _2194;
    wire [3:0] _2197;
    wire [3:0] _2200;
    wire [3:0] _2203;
    wire [3:0] _2206;
    wire _2208;
    wire _2209;
    wire _3446;
    wire _3447;
    wire _3448;
    wire _3449;
    wire _170;
    reg _1879;
    wire [3:0] _2454;
    wire [3:0] _2451;
    wire [3:0] _2448;
    wire [3:0] _2444;
    wire [3:0] _2449;
    wire [3:0] _2452;
    wire [3:0] _2455;
    wire [3:0] _2458;
    wire _2460;
    wire _2461;
    wire _3450;
    wire _3451;
    wire _3452;
    wire _3453;
    wire _171;
    reg _2165;
    wire [3:0] _2739;
    wire [3:0] _2736;
    wire [3:0] _2733;
    wire [3:0] _2730;
    wire [3:0] _2726;
    wire [3:0] _2731;
    wire [3:0] _2734;
    wire [3:0] _2737;
    wire [3:0] _2740;
    wire _2742;
    wire _2743;
    wire _3454;
    wire _3455;
    wire _3456;
    wire _3457;
    wire _172;
    reg _2447;
    wire [3:0] _2472;
    wire [3:0] _2469;
    wire [3:0] _2467;
    wire [3:0] _2470;
    wire [3:0] _2473;
    wire [3:0] _2476;
    wire [3:0] _2479;
    wire [3:0] _2482;
    wire [3:0] _2485;
    wire [3:0] _2488;
    wire _2490;
    wire _2491;
    wire _3458;
    wire _3459;
    wire _3460;
    wire _3461;
    wire _173;
    reg _2161;
    wire [3:0] _2508;
    wire [3:0] _2505;
    wire [3:0] _2502;
    wire [3:0] _2499;
    wire [3:0] _2497;
    wire [3:0] _2500;
    wire [3:0] _2503;
    wire [3:0] _2506;
    wire [3:0] _2509;
    wire [3:0] _2512;
    wire [3:0] _2515;
    wire [3:0] _2518;
    wire _2520;
    wire _2521;
    wire _3462;
    wire _3463;
    wire _3464;
    wire _3465;
    wire _174;
    reg _2184;
    wire [3:0] _2538;
    wire [3:0] _2535;
    wire [3:0] _2532;
    wire [3:0] _2529;
    wire [3:0] _2527;
    wire [3:0] _2530;
    wire [3:0] _2533;
    wire [3:0] _2536;
    wire [3:0] _2539;
    wire [3:0] _2542;
    wire [3:0] _2545;
    wire [3:0] _2548;
    wire _2550;
    wire _2551;
    wire _3466;
    wire _3467;
    wire _3468;
    wire _3469;
    wire _175;
    reg _2214;
    wire [3:0] _2568;
    wire [3:0] _2565;
    wire [3:0] _2562;
    wire [3:0] _2559;
    wire [3:0] _2557;
    wire [3:0] _2560;
    wire [3:0] _2563;
    wire [3:0] _2566;
    wire [3:0] _2569;
    wire [3:0] _2572;
    wire [3:0] _2575;
    wire [3:0] _2578;
    wire _2580;
    wire _2581;
    wire _3470;
    wire _3471;
    wire _3472;
    wire _3473;
    wire _176;
    reg _2244;
    wire [3:0] _2598;
    wire [3:0] _2595;
    wire [3:0] _2592;
    wire [3:0] _2589;
    wire [3:0] _2587;
    wire [3:0] _2590;
    wire [3:0] _2593;
    wire [3:0] _2596;
    wire [3:0] _2599;
    wire [3:0] _2602;
    wire [3:0] _2605;
    wire [3:0] _2608;
    wire _2610;
    wire _2611;
    wire _3474;
    wire _3475;
    wire _3476;
    wire _3477;
    wire _177;
    reg _2274;
    wire [3:0] _2628;
    wire [3:0] _2625;
    wire [3:0] _2622;
    wire [3:0] _2619;
    wire [3:0] _2617;
    wire [3:0] _2620;
    wire [3:0] _2623;
    wire [3:0] _2626;
    wire [3:0] _2629;
    wire [3:0] _2632;
    wire [3:0] _2635;
    wire [3:0] _2638;
    wire _2640;
    wire _2641;
    wire _3478;
    wire _3479;
    wire _3480;
    wire _3481;
    wire _178;
    reg _2304;
    wire [3:0] _2658;
    wire [3:0] _2655;
    wire [3:0] _2652;
    wire [3:0] _2649;
    wire [3:0] _2647;
    wire [3:0] _2650;
    wire [3:0] _2653;
    wire [3:0] _2656;
    wire [3:0] _2659;
    wire [3:0] _2662;
    wire [3:0] _2665;
    wire [3:0] _2668;
    wire _2670;
    wire _2671;
    wire _3482;
    wire _3483;
    wire _3484;
    wire _3485;
    wire _179;
    reg _2334;
    wire [3:0] _2688;
    wire [3:0] _2685;
    wire [3:0] _2682;
    wire [3:0] _2679;
    wire [3:0] _2677;
    wire [3:0] _2680;
    wire [3:0] _2683;
    wire [3:0] _2686;
    wire [3:0] _2689;
    wire [3:0] _2692;
    wire [3:0] _2695;
    wire [3:0] _2698;
    wire _2700;
    wire _2701;
    wire _3486;
    wire _3487;
    wire _3488;
    wire _3489;
    wire _180;
    reg _2364;
    wire [3:0] _2710;
    wire [3:0] _2707;
    wire [3:0] _2705;
    wire [3:0] _2708;
    wire [3:0] _2711;
    wire [3:0] _2714;
    wire [3:0] _2717;
    wire _2719;
    wire _2720;
    wire _3490;
    wire _3491;
    wire _3492;
    wire _3493;
    wire _181;
    reg _2394;
    wire [3:0] _2995;
    wire [3:0] _2992;
    wire [3:0] _2989;
    wire [3:0] _2987;
    wire [3:0] _2990;
    wire [3:0] _2993;
    wire [3:0] _2996;
    wire [3:0] _2999;
    wire _3001;
    wire _3002;
    wire _3494;
    wire _3495;
    wire _3496;
    wire _3497;
    wire _182;
    reg _2676;
    wire [3:0] _2967;
    wire [3:0] _2964;
    wire [3:0] _2961;
    wire [3:0] _2959;
    wire [3:0] _2962;
    wire [3:0] _2965;
    wire [3:0] _2968;
    wire [3:0] _2971;
    wire [3:0] _2974;
    wire [3:0] _2977;
    wire [3:0] _2980;
    wire _2982;
    wire _2983;
    wire _3498;
    wire _3499;
    wire _3500;
    wire _3501;
    wire _183;
    reg _2646;
    wire [3:0] _2937;
    wire [3:0] _2934;
    wire [3:0] _2931;
    wire [3:0] _2929;
    wire [3:0] _2932;
    wire [3:0] _2935;
    wire [3:0] _2938;
    wire [3:0] _2941;
    wire [3:0] _2944;
    wire [3:0] _2947;
    wire [3:0] _2950;
    wire _2952;
    wire _2953;
    wire _3502;
    wire _3503;
    wire _3504;
    wire _3505;
    wire _184;
    reg _2616;
    wire [3:0] _2907;
    wire [3:0] _2904;
    wire [3:0] _2901;
    wire [3:0] _2899;
    wire [3:0] _2902;
    wire [3:0] _2905;
    wire [3:0] _2908;
    wire [3:0] _2911;
    wire [3:0] _2914;
    wire [3:0] _2917;
    wire [3:0] _2920;
    wire _2922;
    wire _2923;
    wire _3506;
    wire _3507;
    wire _3508;
    wire _3509;
    wire _185;
    reg _2586;
    wire [3:0] _2877;
    wire [3:0] _2874;
    wire [3:0] _2871;
    wire [3:0] _2869;
    wire [3:0] _2872;
    wire [3:0] _2875;
    wire [3:0] _2878;
    wire [3:0] _2881;
    wire [3:0] _2884;
    wire [3:0] _2887;
    wire [3:0] _2890;
    wire _2892;
    wire _2893;
    wire _3510;
    wire _3511;
    wire _3512;
    wire _3513;
    wire _186;
    reg _2556;
    wire [3:0] _2847;
    wire [3:0] _2844;
    wire [3:0] _2841;
    wire [3:0] _2839;
    wire [3:0] _2842;
    wire [3:0] _2845;
    wire [3:0] _2848;
    wire [3:0] _2851;
    wire [3:0] _2854;
    wire [3:0] _2857;
    wire [3:0] _2860;
    wire _2862;
    wire _2863;
    wire _3514;
    wire _3515;
    wire _3516;
    wire _3517;
    wire _187;
    reg _2526;
    wire [3:0] _2817;
    wire [3:0] _2814;
    wire [3:0] _2811;
    wire [3:0] _2809;
    wire [3:0] _2812;
    wire [3:0] _2815;
    wire [3:0] _2818;
    wire [3:0] _2821;
    wire [3:0] _2824;
    wire [3:0] _2827;
    wire [3:0] _2830;
    wire _2832;
    wire _2833;
    wire _3518;
    wire _3519;
    wire _3520;
    wire _3521;
    wire _188;
    reg _2496;
    wire [3:0] _2787;
    wire [3:0] _2784;
    wire [3:0] _2781;
    wire [3:0] _2779;
    wire [3:0] _2782;
    wire [3:0] _2785;
    wire [3:0] _2788;
    wire [3:0] _2791;
    wire [3:0] _2794;
    wire [3:0] _2797;
    wire [3:0] _2800;
    wire _2802;
    wire _2803;
    wire _3522;
    wire _3523;
    wire _3524;
    wire _3525;
    wire _189;
    reg _2466;
    wire [3:0] _2757;
    wire [3:0] _2754;
    wire [3:0] _2751;
    wire [3:0] _2749;
    wire [3:0] _2752;
    wire [3:0] _2755;
    wire [3:0] _2758;
    wire [3:0] _2761;
    wire [3:0] _2764;
    wire [3:0] _2767;
    wire [3:0] _2770;
    wire _2772;
    wire _2773;
    wire _3526;
    wire _3527;
    wire _3528;
    wire _3529;
    wire _190;
    reg _2443;
    wire [3:0] _3008;
    wire [3:0] _3006;
    wire [3:0] _3009;
    wire [3:0] _3012;
    wire _3014;
    wire _3015;
    wire _3530;
    wire _3531;
    wire _3532;
    wire _3533;
    wire _191;
    reg _2729;
    wire [3:0] _3021;
    wire [3:0] _3019;
    wire [3:0] _3022;
    wire [3:0] _3025;
    wire [3:0] _3028;
    wire [3:0] _3031;
    wire _3033;
    wire _3034;
    wire _3534;
    wire _3535;
    wire _3536;
    wire _3537;
    wire _192;
    reg _2725;
    wire [3:0] _3040;
    wire [3:0] _3038;
    wire [3:0] _3041;
    wire [3:0] _3044;
    wire [3:0] _3047;
    wire [3:0] _3050;
    wire _3052;
    wire _3053;
    wire _3538;
    wire _3539;
    wire _3540;
    wire _3541;
    wire _193;
    reg _2748;
    wire [3:0] _3059;
    wire [3:0] _3057;
    wire [3:0] _3060;
    wire [3:0] _3063;
    wire [3:0] _3066;
    wire [3:0] _3069;
    wire _3071;
    wire _3072;
    wire _3542;
    wire _3543;
    wire _3544;
    wire _3545;
    wire _194;
    reg _2778;
    wire [3:0] _3078;
    wire [3:0] _3076;
    wire [3:0] _3079;
    wire [3:0] _3082;
    wire [3:0] _3085;
    wire [3:0] _3088;
    wire _3090;
    wire _3091;
    wire _3546;
    wire _3547;
    wire _3548;
    wire _3549;
    wire _195;
    reg _2808;
    wire [3:0] _3097;
    wire [3:0] _3095;
    wire [3:0] _3098;
    wire [3:0] _3101;
    wire [3:0] _3104;
    wire [3:0] _3107;
    wire _3109;
    wire _3110;
    wire _3550;
    wire _3551;
    wire _3552;
    wire _3553;
    wire _196;
    reg _2838;
    wire [3:0] _3116;
    wire [3:0] _3114;
    wire [3:0] _3117;
    wire [3:0] _3120;
    wire [3:0] _3123;
    wire [3:0] _3126;
    wire _3128;
    wire _3129;
    wire _3554;
    wire _3555;
    wire _3556;
    wire _3557;
    wire _197;
    reg _2868;
    wire [3:0] _3135;
    wire [3:0] _3133;
    wire [3:0] _3136;
    wire [3:0] _3139;
    wire [3:0] _3142;
    wire [3:0] _3145;
    wire _3147;
    wire _3148;
    wire _3558;
    wire _3559;
    wire _3560;
    wire _3561;
    wire _198;
    reg _2898;
    wire [3:0] _3154;
    wire [3:0] _3152;
    wire [3:0] _3155;
    wire [3:0] _3158;
    wire [3:0] _3161;
    wire [3:0] _3164;
    wire _3166;
    wire _3167;
    wire _3562;
    wire _3563;
    wire _3564;
    wire _3565;
    wire _199;
    reg _2928;
    wire [3:0] _3567;
    wire [3:0] _3570;
    wire [3:0] _3573;
    wire _3575;
    wire _220;
    wire _221;
    wire _3580;
    wire _3577;
    wire _3578;
    wire _3579;
    wire _3581;
    wire _200;
    reg _2958;
    wire _3576;
    wire gnd;
    wire _3582;
    wire [3:0] _527;
    wire _528;
    wire _529;
    wire _3583;
    wire _201;
    wire [15:0] _227;
    wire [15:0] _230;
    wire [15:0] _233;
    wire [15:0] _236;
    wire [15:0] _239;
    wire [15:0] _242;
    wire [15:0] _245;
    wire [15:0] _248;
    wire [15:0] _251;
    wire [15:0] _254;
    wire [15:0] _257;
    wire [15:0] _260;
    wire [15:0] _263;
    wire [15:0] _266;
    wire [15:0] _269;
    wire [15:0] _272;
    wire [15:0] _275;
    wire [15:0] _278;
    wire [15:0] _281;
    wire [15:0] _284;
    wire [15:0] _287;
    wire [15:0] _290;
    wire [15:0] _293;
    wire [15:0] _296;
    wire [15:0] _299;
    wire [15:0] _302;
    wire [15:0] _305;
    wire [15:0] _308;
    wire [15:0] _311;
    wire [15:0] _314;
    wire [15:0] _317;
    wire [15:0] _320;
    wire [15:0] _323;
    wire [15:0] _326;
    wire [15:0] _329;
    wire [15:0] _332;
    wire [15:0] _335;
    wire [15:0] _338;
    wire [15:0] _341;
    wire [15:0] _344;
    wire [15:0] _347;
    wire [15:0] _350;
    wire [15:0] _353;
    wire [15:0] _356;
    wire [15:0] _359;
    wire [15:0] _362;
    wire [15:0] _365;
    wire [15:0] _368;
    wire [15:0] _371;
    wire [15:0] _374;
    wire [15:0] _377;
    wire [15:0] _380;
    wire [15:0] _383;
    wire [15:0] _386;
    wire [15:0] _389;
    wire [15:0] _392;
    wire [15:0] _395;
    wire [15:0] _398;
    wire [15:0] _401;
    wire [15:0] _404;
    wire [15:0] _407;
    wire [15:0] _410;
    wire [15:0] _413;
    wire [15:0] _416;
    wire [15:0] _419;
    wire [15:0] _422;
    wire [15:0] _425;
    wire [15:0] _428;
    wire [15:0] _431;
    wire [15:0] _434;
    wire [15:0] _437;
    wire [15:0] _440;
    wire [15:0] _443;
    wire [15:0] _446;
    wire [15:0] _449;
    wire [15:0] _452;
    wire [15:0] _455;
    wire [15:0] _458;
    wire [15:0] _461;
    wire [15:0] _464;
    wire [15:0] _467;
    wire [15:0] _470;
    wire [15:0] _473;
    wire [15:0] _476;
    wire [15:0] _479;
    wire [15:0] _482;
    wire [15:0] _485;
    wire [15:0] _488;
    wire [15:0] _491;
    wire [15:0] _494;
    wire [15:0] _497;
    wire [15:0] _500;
    wire [15:0] _503;
    wire [15:0] _506;
    wire [15:0] _509;
    wire [15:0] _512;
    wire [15:0] _515;
    wire [15:0] _518;
    wire [15:0] _521;
    wire [15:0] _524;
    wire _3587;
    wire _219;
    wire _3588;
    wire [30:0] _3585;
    wire [31:0] _3589;
    wire [31:0] _3584;
    wire [3:0] _215;
    wire _216;
    wire _203;
    wire _217;
    wire _205;
    wire _207;
    wire [31:0] _209;
    wire [31:0] _210;
    reg [31:0] _218;
    wire [3:0] _212;
    reg [31:0] _3893;
    assign _3889 = 15'b000000000000000;
    assign _3890 = { _3889,
                     _532 };
    assign _3887 = { _3889,
                     _544 };
    assign _3884 = { _3889,
                     _564 };
    assign _3881 = { _3889,
                     _587 };
    assign _3878 = { _3889,
                     _610 };
    assign _3875 = { _3889,
                     _633 };
    assign _3872 = { _3889,
                     _656 };
    assign _3869 = { _3889,
                     _679 };
    assign _3866 = { _3889,
                     _702 };
    assign _3863 = { _3889,
                     _725 };
    assign _3860 = { _3889,
                     _539 };
    assign _3857 = { _3889,
                     _535 };
    assign _3854 = { _3889,
                     _554 };
    assign _3851 = { _3889,
                     _577 };
    assign _3848 = { _3889,
                     _600 };
    assign _3845 = { _3889,
                     _623 };
    assign _3842 = { _3889,
                     _646 };
    assign _3839 = { _3889,
                     _669 };
    assign _3836 = { _3889,
                     _692 };
    assign _3833 = { _3889,
                     _715 };
    assign _3830 = { _3889,
                     _755 };
    assign _3827 = { _3889,
                     _751 };
    assign _3824 = { _3889,
                     _774 };
    assign _3821 = { _3889,
                     _804 };
    assign _3818 = { _3889,
                     _834 };
    assign _3815 = { _3889,
                     _864 };
    assign _3812 = { _3889,
                     _894 };
    assign _3809 = { _3889,
                     _924 };
    assign _3806 = { _3889,
                     _954 };
    assign _3803 = { _3889,
                     _984 };
    assign _3800 = { _3889,
                     _1037 };
    assign _3797 = { _3889,
                     _1033 };
    assign _3794 = { _3889,
                     _1056 };
    assign _3791 = { _3889,
                     _1086 };
    assign _3788 = { _3889,
                     _1116 };
    assign _3785 = { _3889,
                     _1146 };
    assign _3782 = { _3889,
                     _1176 };
    assign _3779 = { _3889,
                     _1206 };
    assign _3776 = { _3889,
                     _1236 };
    assign _3773 = { _3889,
                     _1266 };
    assign _3770 = { _3889,
                     _1319 };
    assign _3767 = { _3889,
                     _1315 };
    assign _3764 = { _3889,
                     _1338 };
    assign _3761 = { _3889,
                     _1368 };
    assign _3758 = { _3889,
                     _1398 };
    assign _3755 = { _3889,
                     _1428 };
    assign _3752 = { _3889,
                     _1458 };
    assign _3749 = { _3889,
                     _1488 };
    assign _3746 = { _3889,
                     _1518 };
    assign _3743 = { _3889,
                     _1548 };
    assign _3740 = { _3889,
                     _1601 };
    assign _3737 = { _3889,
                     _1597 };
    assign _3734 = { _3889,
                     _1620 };
    assign _3731 = { _3889,
                     _1650 };
    assign _3728 = { _3889,
                     _1680 };
    assign _3725 = { _3889,
                     _1710 };
    assign _3722 = { _3889,
                     _1740 };
    assign _3719 = { _3889,
                     _1770 };
    assign _3716 = { _3889,
                     _1800 };
    assign _3713 = { _3889,
                     _1830 };
    assign _3710 = { _3889,
                     _1883 };
    assign _3707 = { _3889,
                     _1879 };
    assign _3704 = { _3889,
                     _1902 };
    assign _3701 = { _3889,
                     _1932 };
    assign _3698 = { _3889,
                     _1962 };
    assign _3695 = { _3889,
                     _1992 };
    assign _3692 = { _3889,
                     _2022 };
    assign _3689 = { _3889,
                     _2052 };
    assign _3686 = { _3889,
                     _2082 };
    assign _3683 = { _3889,
                     _2112 };
    assign _3680 = { _3889,
                     _2165 };
    assign _3677 = { _3889,
                     _2161 };
    assign _3674 = { _3889,
                     _2184 };
    assign _3671 = { _3889,
                     _2214 };
    assign _3668 = { _3889,
                     _2244 };
    assign _3665 = { _3889,
                     _2274 };
    assign _3662 = { _3889,
                     _2304 };
    assign _3659 = { _3889,
                     _2334 };
    assign _3656 = { _3889,
                     _2364 };
    assign _3653 = { _3889,
                     _2394 };
    assign _3650 = { _3889,
                     _2447 };
    assign _3647 = { _3889,
                     _2443 };
    assign _3644 = { _3889,
                     _2466 };
    assign _3641 = { _3889,
                     _2496 };
    assign _3638 = { _3889,
                     _2526 };
    assign _3635 = { _3889,
                     _2556 };
    assign _3632 = { _3889,
                     _2586 };
    assign _3629 = { _3889,
                     _2616 };
    assign _3626 = { _3889,
                     _2646 };
    assign _3623 = { _3889,
                     _2676 };
    assign _3620 = { _3889,
                     _2729 };
    assign _3617 = { _3889,
                     _2725 };
    assign _3614 = { _3889,
                     _2748 };
    assign _3611 = { _3889,
                     _2778 };
    assign _3608 = { _3889,
                     _2808 };
    assign _3605 = { _3889,
                     _2838 };
    assign _3602 = { _3889,
                     _2868 };
    assign _3599 = { _3889,
                     _2898 };
    assign _3596 = { _3889,
                     _2928 };
    assign _3594 = { _3889,
                     _2958 };
    assign _3597 = _3594 + _3596;
    assign _3600 = _3597 + _3599;
    assign _3603 = _3600 + _3602;
    assign _3606 = _3603 + _3605;
    assign _3609 = _3606 + _3608;
    assign _3612 = _3609 + _3611;
    assign _3615 = _3612 + _3614;
    assign _3618 = _3615 + _3617;
    assign _3621 = _3618 + _3620;
    assign _3624 = _3621 + _3623;
    assign _3627 = _3624 + _3626;
    assign _3630 = _3627 + _3629;
    assign _3633 = _3630 + _3632;
    assign _3636 = _3633 + _3635;
    assign _3639 = _3636 + _3638;
    assign _3642 = _3639 + _3641;
    assign _3645 = _3642 + _3644;
    assign _3648 = _3645 + _3647;
    assign _3651 = _3648 + _3650;
    assign _3654 = _3651 + _3653;
    assign _3657 = _3654 + _3656;
    assign _3660 = _3657 + _3659;
    assign _3663 = _3660 + _3662;
    assign _3666 = _3663 + _3665;
    assign _3669 = _3666 + _3668;
    assign _3672 = _3669 + _3671;
    assign _3675 = _3672 + _3674;
    assign _3678 = _3675 + _3677;
    assign _3681 = _3678 + _3680;
    assign _3684 = _3681 + _3683;
    assign _3687 = _3684 + _3686;
    assign _3690 = _3687 + _3689;
    assign _3693 = _3690 + _3692;
    assign _3696 = _3693 + _3695;
    assign _3699 = _3696 + _3698;
    assign _3702 = _3699 + _3701;
    assign _3705 = _3702 + _3704;
    assign _3708 = _3705 + _3707;
    assign _3711 = _3708 + _3710;
    assign _3714 = _3711 + _3713;
    assign _3717 = _3714 + _3716;
    assign _3720 = _3717 + _3719;
    assign _3723 = _3720 + _3722;
    assign _3726 = _3723 + _3725;
    assign _3729 = _3726 + _3728;
    assign _3732 = _3729 + _3731;
    assign _3735 = _3732 + _3734;
    assign _3738 = _3735 + _3737;
    assign _3741 = _3738 + _3740;
    assign _3744 = _3741 + _3743;
    assign _3747 = _3744 + _3746;
    assign _3750 = _3747 + _3749;
    assign _3753 = _3750 + _3752;
    assign _3756 = _3753 + _3755;
    assign _3759 = _3756 + _3758;
    assign _3762 = _3759 + _3761;
    assign _3765 = _3762 + _3764;
    assign _3768 = _3765 + _3767;
    assign _3771 = _3768 + _3770;
    assign _3774 = _3771 + _3773;
    assign _3777 = _3774 + _3776;
    assign _3780 = _3777 + _3779;
    assign _3783 = _3780 + _3782;
    assign _3786 = _3783 + _3785;
    assign _3789 = _3786 + _3788;
    assign _3792 = _3789 + _3791;
    assign _3795 = _3792 + _3794;
    assign _3798 = _3795 + _3797;
    assign _3801 = _3798 + _3800;
    assign _3804 = _3801 + _3803;
    assign _3807 = _3804 + _3806;
    assign _3810 = _3807 + _3809;
    assign _3813 = _3810 + _3812;
    assign _3816 = _3813 + _3815;
    assign _3819 = _3816 + _3818;
    assign _3822 = _3819 + _3821;
    assign _3825 = _3822 + _3824;
    assign _3828 = _3825 + _3827;
    assign _3831 = _3828 + _3830;
    assign _3834 = _3831 + _3833;
    assign _3837 = _3834 + _3836;
    assign _3840 = _3837 + _3839;
    assign _3843 = _3840 + _3842;
    assign _3846 = _3843 + _3845;
    assign _3849 = _3846 + _3848;
    assign _3852 = _3849 + _3851;
    assign _3855 = _3852 + _3854;
    assign _3858 = _3855 + _3857;
    assign _3861 = _3858 + _3860;
    assign _3864 = _3861 + _3863;
    assign _3867 = _3864 + _3866;
    assign _3870 = _3867 + _3869;
    assign _3873 = _3870 + _3872;
    assign _3876 = _3873 + _3875;
    assign _3879 = _3876 + _3878;
    assign _3882 = _3879 + _3881;
    assign _3885 = _3882 + _3884;
    assign _3888 = _3885 + _3887;
    assign _3891 = _3888 + _3890;
    assign _3592 = 16'b0000000000000000;
    assign _3892 = { _3592,
                     _3891 };
    assign _525 = _223 + _524;
    assign _225 = _221 ? _3592 : _223;
    assign _526 = _219 ? _525 : _225;
    assign _1 = _526;
    always @(posedge _207) begin
        if (_221)
            _223 <= _3592;
        else
            _223 <= _1;
    end
    assign _3591 = { _3592,
                     _223 };
    assign _550 = _219 ? _549 : gnd;
    assign _551 = _529 ? gnd : _550;
    assign _2 = _551;
    assign _523 = { _3889,
                    _2 };
    assign _573 = _219 ? _572 : gnd;
    assign _574 = _529 ? gnd : _573;
    assign _3 = _574;
    assign _520 = { _3889,
                    _3 };
    assign _596 = _219 ? _595 : gnd;
    assign _597 = _529 ? gnd : _596;
    assign _4 = _597;
    assign _517 = { _3889,
                    _4 };
    assign _619 = _219 ? _618 : gnd;
    assign _620 = _529 ? gnd : _619;
    assign _5 = _620;
    assign _514 = { _3889,
                    _5 };
    assign _642 = _219 ? _641 : gnd;
    assign _643 = _529 ? gnd : _642;
    assign _6 = _643;
    assign _511 = { _3889,
                    _6 };
    assign _665 = _219 ? _664 : gnd;
    assign _666 = _529 ? gnd : _665;
    assign _7 = _666;
    assign _508 = { _3889,
                    _7 };
    assign _688 = _219 ? _687 : gnd;
    assign _689 = _529 ? gnd : _688;
    assign _8 = _689;
    assign _505 = { _3889,
                    _8 };
    assign _711 = _219 ? _710 : gnd;
    assign _712 = _529 ? gnd : _711;
    assign _9 = _712;
    assign _502 = { _3889,
                    _9 };
    assign _734 = _219 ? _733 : gnd;
    assign _735 = _529 ? gnd : _734;
    assign _10 = _735;
    assign _499 = { _3889,
                    _10 };
    assign _747 = _219 ? _746 : gnd;
    assign _748 = _529 ? gnd : _747;
    assign _11 = _748;
    assign _496 = { _3889,
                    _11 };
    assign _770 = _219 ? _769 : gnd;
    assign _771 = _529 ? gnd : _770;
    assign _12 = _771;
    assign _493 = { _3889,
                    _12 };
    assign _800 = _219 ? _799 : gnd;
    assign _801 = _529 ? gnd : _800;
    assign _13 = _801;
    assign _490 = { _3889,
                    _13 };
    assign _830 = _219 ? _829 : gnd;
    assign _831 = _529 ? gnd : _830;
    assign _14 = _831;
    assign _487 = { _3889,
                    _14 };
    assign _860 = _219 ? _859 : gnd;
    assign _861 = _529 ? gnd : _860;
    assign _15 = _861;
    assign _484 = { _3889,
                    _15 };
    assign _890 = _219 ? _889 : gnd;
    assign _891 = _529 ? gnd : _890;
    assign _16 = _891;
    assign _481 = { _3889,
                    _16 };
    assign _920 = _219 ? _919 : gnd;
    assign _921 = _529 ? gnd : _920;
    assign _17 = _921;
    assign _478 = { _3889,
                    _17 };
    assign _950 = _219 ? _949 : gnd;
    assign _951 = _529 ? gnd : _950;
    assign _18 = _951;
    assign _475 = { _3889,
                    _18 };
    assign _980 = _219 ? _979 : gnd;
    assign _981 = _529 ? gnd : _980;
    assign _19 = _981;
    assign _472 = { _3889,
                    _19 };
    assign _1010 = _219 ? _1009 : gnd;
    assign _1011 = _529 ? gnd : _1010;
    assign _20 = _1011;
    assign _469 = { _3889,
                    _20 };
    assign _1029 = _219 ? _1028 : gnd;
    assign _1030 = _529 ? gnd : _1029;
    assign _21 = _1030;
    assign _466 = { _3889,
                    _21 };
    assign _1052 = _219 ? _1051 : gnd;
    assign _1053 = _529 ? gnd : _1052;
    assign _22 = _1053;
    assign _463 = { _3889,
                    _22 };
    assign _1082 = _219 ? _1081 : gnd;
    assign _1083 = _529 ? gnd : _1082;
    assign _23 = _1083;
    assign _460 = { _3889,
                    _23 };
    assign _1112 = _219 ? _1111 : gnd;
    assign _1113 = _529 ? gnd : _1112;
    assign _24 = _1113;
    assign _457 = { _3889,
                    _24 };
    assign _1142 = _219 ? _1141 : gnd;
    assign _1143 = _529 ? gnd : _1142;
    assign _25 = _1143;
    assign _454 = { _3889,
                    _25 };
    assign _1172 = _219 ? _1171 : gnd;
    assign _1173 = _529 ? gnd : _1172;
    assign _26 = _1173;
    assign _451 = { _3889,
                    _26 };
    assign _1202 = _219 ? _1201 : gnd;
    assign _1203 = _529 ? gnd : _1202;
    assign _27 = _1203;
    assign _448 = { _3889,
                    _27 };
    assign _1232 = _219 ? _1231 : gnd;
    assign _1233 = _529 ? gnd : _1232;
    assign _28 = _1233;
    assign _445 = { _3889,
                    _28 };
    assign _1262 = _219 ? _1261 : gnd;
    assign _1263 = _529 ? gnd : _1262;
    assign _29 = _1263;
    assign _442 = { _3889,
                    _29 };
    assign _1292 = _219 ? _1291 : gnd;
    assign _1293 = _529 ? gnd : _1292;
    assign _30 = _1293;
    assign _439 = { _3889,
                    _30 };
    assign _1311 = _219 ? _1310 : gnd;
    assign _1312 = _529 ? gnd : _1311;
    assign _31 = _1312;
    assign _436 = { _3889,
                    _31 };
    assign _1334 = _219 ? _1333 : gnd;
    assign _1335 = _529 ? gnd : _1334;
    assign _32 = _1335;
    assign _433 = { _3889,
                    _32 };
    assign _1364 = _219 ? _1363 : gnd;
    assign _1365 = _529 ? gnd : _1364;
    assign _33 = _1365;
    assign _430 = { _3889,
                    _33 };
    assign _1394 = _219 ? _1393 : gnd;
    assign _1395 = _529 ? gnd : _1394;
    assign _34 = _1395;
    assign _427 = { _3889,
                    _34 };
    assign _1424 = _219 ? _1423 : gnd;
    assign _1425 = _529 ? gnd : _1424;
    assign _35 = _1425;
    assign _424 = { _3889,
                    _35 };
    assign _1454 = _219 ? _1453 : gnd;
    assign _1455 = _529 ? gnd : _1454;
    assign _36 = _1455;
    assign _421 = { _3889,
                    _36 };
    assign _1484 = _219 ? _1483 : gnd;
    assign _1485 = _529 ? gnd : _1484;
    assign _37 = _1485;
    assign _418 = { _3889,
                    _37 };
    assign _1514 = _219 ? _1513 : gnd;
    assign _1515 = _529 ? gnd : _1514;
    assign _38 = _1515;
    assign _415 = { _3889,
                    _38 };
    assign _1544 = _219 ? _1543 : gnd;
    assign _1545 = _529 ? gnd : _1544;
    assign _39 = _1545;
    assign _412 = { _3889,
                    _39 };
    assign _1574 = _219 ? _1573 : gnd;
    assign _1575 = _529 ? gnd : _1574;
    assign _40 = _1575;
    assign _409 = { _3889,
                    _40 };
    assign _1593 = _219 ? _1592 : gnd;
    assign _1594 = _529 ? gnd : _1593;
    assign _41 = _1594;
    assign _406 = { _3889,
                    _41 };
    assign _1616 = _219 ? _1615 : gnd;
    assign _1617 = _529 ? gnd : _1616;
    assign _42 = _1617;
    assign _403 = { _3889,
                    _42 };
    assign _1646 = _219 ? _1645 : gnd;
    assign _1647 = _529 ? gnd : _1646;
    assign _43 = _1647;
    assign _400 = { _3889,
                    _43 };
    assign _1676 = _219 ? _1675 : gnd;
    assign _1677 = _529 ? gnd : _1676;
    assign _44 = _1677;
    assign _397 = { _3889,
                    _44 };
    assign _1706 = _219 ? _1705 : gnd;
    assign _1707 = _529 ? gnd : _1706;
    assign _45 = _1707;
    assign _394 = { _3889,
                    _45 };
    assign _1736 = _219 ? _1735 : gnd;
    assign _1737 = _529 ? gnd : _1736;
    assign _46 = _1737;
    assign _391 = { _3889,
                    _46 };
    assign _1766 = _219 ? _1765 : gnd;
    assign _1767 = _529 ? gnd : _1766;
    assign _47 = _1767;
    assign _388 = { _3889,
                    _47 };
    assign _1796 = _219 ? _1795 : gnd;
    assign _1797 = _529 ? gnd : _1796;
    assign _48 = _1797;
    assign _385 = { _3889,
                    _48 };
    assign _1826 = _219 ? _1825 : gnd;
    assign _1827 = _529 ? gnd : _1826;
    assign _49 = _1827;
    assign _382 = { _3889,
                    _49 };
    assign _1856 = _219 ? _1855 : gnd;
    assign _1857 = _529 ? gnd : _1856;
    assign _50 = _1857;
    assign _379 = { _3889,
                    _50 };
    assign _1875 = _219 ? _1874 : gnd;
    assign _1876 = _529 ? gnd : _1875;
    assign _51 = _1876;
    assign _376 = { _3889,
                    _51 };
    assign _1898 = _219 ? _1897 : gnd;
    assign _1899 = _529 ? gnd : _1898;
    assign _52 = _1899;
    assign _373 = { _3889,
                    _52 };
    assign _1928 = _219 ? _1927 : gnd;
    assign _1929 = _529 ? gnd : _1928;
    assign _53 = _1929;
    assign _370 = { _3889,
                    _53 };
    assign _1958 = _219 ? _1957 : gnd;
    assign _1959 = _529 ? gnd : _1958;
    assign _54 = _1959;
    assign _367 = { _3889,
                    _54 };
    assign _1988 = _219 ? _1987 : gnd;
    assign _1989 = _529 ? gnd : _1988;
    assign _55 = _1989;
    assign _364 = { _3889,
                    _55 };
    assign _2018 = _219 ? _2017 : gnd;
    assign _2019 = _529 ? gnd : _2018;
    assign _56 = _2019;
    assign _361 = { _3889,
                    _56 };
    assign _2048 = _219 ? _2047 : gnd;
    assign _2049 = _529 ? gnd : _2048;
    assign _57 = _2049;
    assign _358 = { _3889,
                    _57 };
    assign _2078 = _219 ? _2077 : gnd;
    assign _2079 = _529 ? gnd : _2078;
    assign _58 = _2079;
    assign _355 = { _3889,
                    _58 };
    assign _2108 = _219 ? _2107 : gnd;
    assign _2109 = _529 ? gnd : _2108;
    assign _59 = _2109;
    assign _352 = { _3889,
                    _59 };
    assign _2138 = _219 ? _2137 : gnd;
    assign _2139 = _529 ? gnd : _2138;
    assign _60 = _2139;
    assign _349 = { _3889,
                    _60 };
    assign _2157 = _219 ? _2156 : gnd;
    assign _2158 = _529 ? gnd : _2157;
    assign _61 = _2158;
    assign _346 = { _3889,
                    _61 };
    assign _2180 = _219 ? _2179 : gnd;
    assign _2181 = _529 ? gnd : _2180;
    assign _62 = _2181;
    assign _343 = { _3889,
                    _62 };
    assign _2210 = _219 ? _2209 : gnd;
    assign _2211 = _529 ? gnd : _2210;
    assign _63 = _2211;
    assign _340 = { _3889,
                    _63 };
    assign _2240 = _219 ? _2239 : gnd;
    assign _2241 = _529 ? gnd : _2240;
    assign _64 = _2241;
    assign _337 = { _3889,
                    _64 };
    assign _2270 = _219 ? _2269 : gnd;
    assign _2271 = _529 ? gnd : _2270;
    assign _65 = _2271;
    assign _334 = { _3889,
                    _65 };
    assign _2300 = _219 ? _2299 : gnd;
    assign _2301 = _529 ? gnd : _2300;
    assign _66 = _2301;
    assign _331 = { _3889,
                    _66 };
    assign _2330 = _219 ? _2329 : gnd;
    assign _2331 = _529 ? gnd : _2330;
    assign _67 = _2331;
    assign _328 = { _3889,
                    _67 };
    assign _2360 = _219 ? _2359 : gnd;
    assign _2361 = _529 ? gnd : _2360;
    assign _68 = _2361;
    assign _325 = { _3889,
                    _68 };
    assign _2390 = _219 ? _2389 : gnd;
    assign _2391 = _529 ? gnd : _2390;
    assign _69 = _2391;
    assign _322 = { _3889,
                    _69 };
    assign _2420 = _219 ? _2419 : gnd;
    assign _2421 = _529 ? gnd : _2420;
    assign _70 = _2421;
    assign _319 = { _3889,
                    _70 };
    assign _2439 = _219 ? _2438 : gnd;
    assign _2440 = _529 ? gnd : _2439;
    assign _71 = _2440;
    assign _316 = { _3889,
                    _71 };
    assign _2462 = _219 ? _2461 : gnd;
    assign _2463 = _529 ? gnd : _2462;
    assign _72 = _2463;
    assign _313 = { _3889,
                    _72 };
    assign _2492 = _219 ? _2491 : gnd;
    assign _2493 = _529 ? gnd : _2492;
    assign _73 = _2493;
    assign _310 = { _3889,
                    _73 };
    assign _2522 = _219 ? _2521 : gnd;
    assign _2523 = _529 ? gnd : _2522;
    assign _74 = _2523;
    assign _307 = { _3889,
                    _74 };
    assign _2552 = _219 ? _2551 : gnd;
    assign _2553 = _529 ? gnd : _2552;
    assign _75 = _2553;
    assign _304 = { _3889,
                    _75 };
    assign _2582 = _219 ? _2581 : gnd;
    assign _2583 = _529 ? gnd : _2582;
    assign _76 = _2583;
    assign _301 = { _3889,
                    _76 };
    assign _2612 = _219 ? _2611 : gnd;
    assign _2613 = _529 ? gnd : _2612;
    assign _77 = _2613;
    assign _298 = { _3889,
                    _77 };
    assign _2642 = _219 ? _2641 : gnd;
    assign _2643 = _529 ? gnd : _2642;
    assign _78 = _2643;
    assign _295 = { _3889,
                    _78 };
    assign _2672 = _219 ? _2671 : gnd;
    assign _2673 = _529 ? gnd : _2672;
    assign _79 = _2673;
    assign _292 = { _3889,
                    _79 };
    assign _2702 = _219 ? _2701 : gnd;
    assign _2703 = _529 ? gnd : _2702;
    assign _80 = _2703;
    assign _289 = { _3889,
                    _80 };
    assign _2721 = _219 ? _2720 : gnd;
    assign _2722 = _529 ? gnd : _2721;
    assign _81 = _2722;
    assign _286 = { _3889,
                    _81 };
    assign _2744 = _219 ? _2743 : gnd;
    assign _2745 = _529 ? gnd : _2744;
    assign _82 = _2745;
    assign _283 = { _3889,
                    _82 };
    assign _2774 = _219 ? _2773 : gnd;
    assign _2775 = _529 ? gnd : _2774;
    assign _83 = _2775;
    assign _280 = { _3889,
                    _83 };
    assign _2804 = _219 ? _2803 : gnd;
    assign _2805 = _529 ? gnd : _2804;
    assign _84 = _2805;
    assign _277 = { _3889,
                    _84 };
    assign _2834 = _219 ? _2833 : gnd;
    assign _2835 = _529 ? gnd : _2834;
    assign _85 = _2835;
    assign _274 = { _3889,
                    _85 };
    assign _2864 = _219 ? _2863 : gnd;
    assign _2865 = _529 ? gnd : _2864;
    assign _86 = _2865;
    assign _271 = { _3889,
                    _86 };
    assign _2894 = _219 ? _2893 : gnd;
    assign _2895 = _529 ? gnd : _2894;
    assign _87 = _2895;
    assign _268 = { _3889,
                    _87 };
    assign _2924 = _219 ? _2923 : gnd;
    assign _2925 = _529 ? gnd : _2924;
    assign _88 = _2925;
    assign _265 = { _3889,
                    _88 };
    assign _2954 = _219 ? _2953 : gnd;
    assign _2955 = _529 ? gnd : _2954;
    assign _89 = _2955;
    assign _262 = { _3889,
                    _89 };
    assign _2984 = _219 ? _2983 : gnd;
    assign _2985 = _529 ? gnd : _2984;
    assign _90 = _2985;
    assign _259 = { _3889,
                    _90 };
    assign _3003 = _219 ? _3002 : gnd;
    assign _3004 = _529 ? gnd : _3003;
    assign _91 = _3004;
    assign _256 = { _3889,
                    _91 };
    assign _3016 = _219 ? _3015 : gnd;
    assign _3017 = _529 ? gnd : _3016;
    assign _92 = _3017;
    assign _253 = { _3889,
                    _92 };
    assign _3035 = _219 ? _3034 : gnd;
    assign _3036 = _529 ? gnd : _3035;
    assign _93 = _3036;
    assign _250 = { _3889,
                    _93 };
    assign _3054 = _219 ? _3053 : gnd;
    assign _3055 = _529 ? gnd : _3054;
    assign _94 = _3055;
    assign _247 = { _3889,
                    _94 };
    assign _3073 = _219 ? _3072 : gnd;
    assign _3074 = _529 ? gnd : _3073;
    assign _95 = _3074;
    assign _244 = { _3889,
                    _95 };
    assign _3092 = _219 ? _3091 : gnd;
    assign _3093 = _529 ? gnd : _3092;
    assign _96 = _3093;
    assign _241 = { _3889,
                    _96 };
    assign _3111 = _219 ? _3110 : gnd;
    assign _3112 = _529 ? gnd : _3111;
    assign _97 = _3112;
    assign _238 = { _3889,
                    _97 };
    assign _3130 = _219 ? _3129 : gnd;
    assign _3131 = _529 ? gnd : _3130;
    assign _98 = _3131;
    assign _235 = { _3889,
                    _98 };
    assign _3149 = _219 ? _3148 : gnd;
    assign _3150 = _529 ? gnd : _3149;
    assign _99 = _3150;
    assign _232 = { _3889,
                    _99 };
    assign _3168 = _219 ? _3167 : gnd;
    assign _3169 = _529 ? gnd : _3168;
    assign _100 = _3169;
    assign _229 = { _3889,
                    _100 };
    assign _3574 = 4'b0100;
    assign _3571 = 3'b000;
    assign _3572 = { _3571,
                     _2646 };
    assign _3569 = { _3571,
                     _2676 };
    assign _2927 = 1'b0;
    assign _3163 = { _3571,
                     _2616 };
    assign _3160 = { _3571,
                     _2646 };
    assign _3157 = { _3571,
                     _2676 };
    assign _3144 = { _3571,
                     _2586 };
    assign _3141 = { _3571,
                     _2616 };
    assign _3138 = { _3571,
                     _2646 };
    assign _3125 = { _3571,
                     _2556 };
    assign _3122 = { _3571,
                     _2586 };
    assign _3119 = { _3571,
                     _2616 };
    assign _3106 = { _3571,
                     _2526 };
    assign _3103 = { _3571,
                     _2556 };
    assign _3100 = { _3571,
                     _2586 };
    assign _3087 = { _3571,
                     _2496 };
    assign _3084 = { _3571,
                     _2526 };
    assign _3081 = { _3571,
                     _2556 };
    assign _3068 = { _3571,
                     _2466 };
    assign _3065 = { _3571,
                     _2496 };
    assign _3062 = { _3571,
                     _2526 };
    assign _3049 = { _3571,
                     _2443 };
    assign _3046 = { _3571,
                     _2466 };
    assign _3043 = { _3571,
                     _2496 };
    assign _3030 = { _3571,
                     _2447 };
    assign _3027 = { _3571,
                     _2443 };
    assign _3024 = { _3571,
                     _2466 };
    assign _3011 = { _3571,
                     _2447 };
    assign _2769 = { _3571,
                     _2165 };
    assign _2766 = { _3571,
                     _2161 };
    assign _2763 = { _3571,
                     _2184 };
    assign _2760 = { _3571,
                     _2447 };
    assign _2799 = { _3571,
                     _2161 };
    assign _2796 = { _3571,
                     _2184 };
    assign _2793 = { _3571,
                     _2214 };
    assign _2790 = { _3571,
                     _2443 };
    assign _2829 = { _3571,
                     _2184 };
    assign _2826 = { _3571,
                     _2214 };
    assign _2823 = { _3571,
                     _2244 };
    assign _2820 = { _3571,
                     _2466 };
    assign _2859 = { _3571,
                     _2214 };
    assign _2856 = { _3571,
                     _2244 };
    assign _2853 = { _3571,
                     _2274 };
    assign _2850 = { _3571,
                     _2496 };
    assign _2889 = { _3571,
                     _2244 };
    assign _2886 = { _3571,
                     _2274 };
    assign _2883 = { _3571,
                     _2304 };
    assign _2880 = { _3571,
                     _2526 };
    assign _2919 = { _3571,
                     _2274 };
    assign _2916 = { _3571,
                     _2304 };
    assign _2913 = { _3571,
                     _2334 };
    assign _2910 = { _3571,
                     _2556 };
    assign _2949 = { _3571,
                     _2304 };
    assign _2946 = { _3571,
                     _2334 };
    assign _2943 = { _3571,
                     _2364 };
    assign _2940 = { _3571,
                     _2586 };
    assign _2979 = { _3571,
                     _2334 };
    assign _2976 = { _3571,
                     _2364 };
    assign _2973 = { _3571,
                     _2394 };
    assign _2970 = { _3571,
                     _2616 };
    assign _2998 = { _3571,
                     _2364 };
    assign _2716 = { _3571,
                     _2082 };
    assign _2713 = { _3571,
                     _2112 };
    assign _2697 = { _3571,
                     _2052 };
    assign _2694 = { _3571,
                     _2082 };
    assign _2691 = { _3571,
                     _2112 };
    assign _2667 = { _3571,
                     _2022 };
    assign _2664 = { _3571,
                     _2052 };
    assign _2661 = { _3571,
                     _2082 };
    assign _2637 = { _3571,
                     _1992 };
    assign _2634 = { _3571,
                     _2022 };
    assign _2631 = { _3571,
                     _2052 };
    assign _2607 = { _3571,
                     _1962 };
    assign _2604 = { _3571,
                     _1992 };
    assign _2601 = { _3571,
                     _2022 };
    assign _2577 = { _3571,
                     _1932 };
    assign _2574 = { _3571,
                     _1962 };
    assign _2571 = { _3571,
                     _1992 };
    assign _2547 = { _3571,
                     _1902 };
    assign _2544 = { _3571,
                     _1932 };
    assign _2541 = { _3571,
                     _1962 };
    assign _2517 = { _3571,
                     _1879 };
    assign _2514 = { _3571,
                     _1902 };
    assign _2511 = { _3571,
                     _1932 };
    assign _2487 = { _3571,
                     _1883 };
    assign _2484 = { _3571,
                     _1879 };
    assign _2481 = { _3571,
                     _1902 };
    assign _2478 = { _3571,
                     _2165 };
    assign _2475 = { _3571,
                     _2184 };
    assign _2457 = { _3571,
                     _1883 };
    assign _2205 = { _3571,
                     _1601 };
    assign _2202 = { _3571,
                     _1597 };
    assign _2199 = { _3571,
                     _1620 };
    assign _2196 = { _3571,
                     _1883 };
    assign _2235 = { _3571,
                     _1597 };
    assign _2232 = { _3571,
                     _1620 };
    assign _2229 = { _3571,
                     _1650 };
    assign _2226 = { _3571,
                     _1879 };
    assign _2265 = { _3571,
                     _1620 };
    assign _2262 = { _3571,
                     _1650 };
    assign _2259 = { _3571,
                     _1680 };
    assign _2256 = { _3571,
                     _1902 };
    assign _2295 = { _3571,
                     _1650 };
    assign _2292 = { _3571,
                     _1680 };
    assign _2289 = { _3571,
                     _1710 };
    assign _2286 = { _3571,
                     _1932 };
    assign _2325 = { _3571,
                     _1680 };
    assign _2322 = { _3571,
                     _1710 };
    assign _2319 = { _3571,
                     _1740 };
    assign _2316 = { _3571,
                     _1962 };
    assign _2355 = { _3571,
                     _1710 };
    assign _2352 = { _3571,
                     _1740 };
    assign _2349 = { _3571,
                     _1770 };
    assign _2346 = { _3571,
                     _1992 };
    assign _2385 = { _3571,
                     _1740 };
    assign _2382 = { _3571,
                     _1770 };
    assign _2379 = { _3571,
                     _1800 };
    assign _2376 = { _3571,
                     _2022 };
    assign _2415 = { _3571,
                     _1770 };
    assign _2412 = { _3571,
                     _1800 };
    assign _2409 = { _3571,
                     _1830 };
    assign _2406 = { _3571,
                     _2052 };
    assign _2434 = { _3571,
                     _1800 };
    assign _2152 = { _3571,
                     _1518 };
    assign _2149 = { _3571,
                     _1548 };
    assign _2133 = { _3571,
                     _1488 };
    assign _2130 = { _3571,
                     _1518 };
    assign _2127 = { _3571,
                     _1548 };
    assign _2103 = { _3571,
                     _1458 };
    assign _2100 = { _3571,
                     _1488 };
    assign _2097 = { _3571,
                     _1518 };
    assign _2073 = { _3571,
                     _1428 };
    assign _2070 = { _3571,
                     _1458 };
    assign _2067 = { _3571,
                     _1488 };
    assign _2043 = { _3571,
                     _1398 };
    assign _2040 = { _3571,
                     _1428 };
    assign _2037 = { _3571,
                     _1458 };
    assign _2013 = { _3571,
                     _1368 };
    assign _2010 = { _3571,
                     _1398 };
    assign _2007 = { _3571,
                     _1428 };
    assign _1983 = { _3571,
                     _1338 };
    assign _1980 = { _3571,
                     _1368 };
    assign _1977 = { _3571,
                     _1398 };
    assign _1953 = { _3571,
                     _1315 };
    assign _1950 = { _3571,
                     _1338 };
    assign _1947 = { _3571,
                     _1368 };
    assign _1923 = { _3571,
                     _1319 };
    assign _1920 = { _3571,
                     _1315 };
    assign _1917 = { _3571,
                     _1338 };
    assign _1914 = { _3571,
                     _1601 };
    assign _1911 = { _3571,
                     _1620 };
    assign _1893 = { _3571,
                     _1319 };
    assign _1641 = { _3571,
                     _1037 };
    assign _1638 = { _3571,
                     _1033 };
    assign _1635 = { _3571,
                     _1056 };
    assign _1632 = { _3571,
                     _1319 };
    assign _1671 = { _3571,
                     _1033 };
    assign _1668 = { _3571,
                     _1056 };
    assign _1665 = { _3571,
                     _1086 };
    assign _1662 = { _3571,
                     _1315 };
    assign _1701 = { _3571,
                     _1056 };
    assign _1698 = { _3571,
                     _1086 };
    assign _1695 = { _3571,
                     _1116 };
    assign _1692 = { _3571,
                     _1338 };
    assign _1731 = { _3571,
                     _1086 };
    assign _1728 = { _3571,
                     _1116 };
    assign _1725 = { _3571,
                     _1146 };
    assign _1722 = { _3571,
                     _1368 };
    assign _1761 = { _3571,
                     _1116 };
    assign _1758 = { _3571,
                     _1146 };
    assign _1755 = { _3571,
                     _1176 };
    assign _1752 = { _3571,
                     _1398 };
    assign _1791 = { _3571,
                     _1146 };
    assign _1788 = { _3571,
                     _1176 };
    assign _1785 = { _3571,
                     _1206 };
    assign _1782 = { _3571,
                     _1428 };
    assign _1821 = { _3571,
                     _1176 };
    assign _1818 = { _3571,
                     _1206 };
    assign _1815 = { _3571,
                     _1236 };
    assign _1812 = { _3571,
                     _1458 };
    assign _1851 = { _3571,
                     _1206 };
    assign _1848 = { _3571,
                     _1236 };
    assign _1845 = { _3571,
                     _1266 };
    assign _1842 = { _3571,
                     _1488 };
    assign _1870 = { _3571,
                     _1236 };
    assign _1588 = { _3571,
                     _954 };
    assign _1585 = { _3571,
                     _984 };
    assign _1569 = { _3571,
                     _924 };
    assign _1566 = { _3571,
                     _954 };
    assign _1563 = { _3571,
                     _984 };
    assign _1539 = { _3571,
                     _894 };
    assign _1536 = { _3571,
                     _924 };
    assign _1533 = { _3571,
                     _954 };
    assign _1509 = { _3571,
                     _864 };
    assign _1506 = { _3571,
                     _894 };
    assign _1503 = { _3571,
                     _924 };
    assign _1479 = { _3571,
                     _834 };
    assign _1476 = { _3571,
                     _864 };
    assign _1473 = { _3571,
                     _894 };
    assign _1449 = { _3571,
                     _804 };
    assign _1446 = { _3571,
                     _834 };
    assign _1443 = { _3571,
                     _864 };
    assign _1419 = { _3571,
                     _774 };
    assign _1416 = { _3571,
                     _804 };
    assign _1413 = { _3571,
                     _834 };
    assign _1389 = { _3571,
                     _751 };
    assign _1386 = { _3571,
                     _774 };
    assign _1383 = { _3571,
                     _804 };
    assign _1359 = { _3571,
                     _755 };
    assign _1356 = { _3571,
                     _751 };
    assign _1353 = { _3571,
                     _774 };
    assign _1350 = { _3571,
                     _1037 };
    assign _1347 = { _3571,
                     _1056 };
    assign _1329 = { _3571,
                     _755 };
    assign _1077 = { _3571,
                     _539 };
    assign _1074 = { _3571,
                     _535 };
    assign _1071 = { _3571,
                     _554 };
    assign _1068 = { _3571,
                     _755 };
    assign _1107 = { _3571,
                     _535 };
    assign _1104 = { _3571,
                     _554 };
    assign _1101 = { _3571,
                     _577 };
    assign _1098 = { _3571,
                     _751 };
    assign _1137 = { _3571,
                     _554 };
    assign _1134 = { _3571,
                     _577 };
    assign _1131 = { _3571,
                     _600 };
    assign _1128 = { _3571,
                     _774 };
    assign _1167 = { _3571,
                     _577 };
    assign _1164 = { _3571,
                     _600 };
    assign _1161 = { _3571,
                     _623 };
    assign _1158 = { _3571,
                     _804 };
    assign _1197 = { _3571,
                     _600 };
    assign _1194 = { _3571,
                     _623 };
    assign _1191 = { _3571,
                     _646 };
    assign _1188 = { _3571,
                     _834 };
    assign _1227 = { _3571,
                     _623 };
    assign _1224 = { _3571,
                     _646 };
    assign _1221 = { _3571,
                     _669 };
    assign _1218 = { _3571,
                     _864 };
    assign _1257 = { _3571,
                     _646 };
    assign _1254 = { _3571,
                     _669 };
    assign _1251 = { _3571,
                     _692 };
    assign _1248 = { _3571,
                     _894 };
    assign _1287 = { _3571,
                     _669 };
    assign _1284 = { _3571,
                     _692 };
    assign _1281 = { _3571,
                     _715 };
    assign _1278 = { _3571,
                     _924 };
    assign _1306 = { _3571,
                     _692 };
    assign _1024 = { _3571,
                     _702 };
    assign _1021 = { _3571,
                     _725 };
    assign _1005 = { _3571,
                     _679 };
    assign _1002 = { _3571,
                     _702 };
    assign _999 = { _3571,
                    _725 };
    assign _975 = { _3571,
                    _656 };
    assign _972 = { _3571,
                    _679 };
    assign _969 = { _3571,
                    _702 };
    assign _945 = { _3571,
                    _633 };
    assign _942 = { _3571,
                    _656 };
    assign _939 = { _3571,
                    _679 };
    assign _915 = { _3571,
                    _610 };
    assign _912 = { _3571,
                    _633 };
    assign _909 = { _3571,
                    _656 };
    assign _885 = { _3571,
                    _587 };
    assign _882 = { _3571,
                    _610 };
    assign _879 = { _3571,
                    _633 };
    assign _855 = { _3571,
                    _564 };
    assign _852 = { _3571,
                    _587 };
    assign _849 = { _3571,
                    _610 };
    assign _825 = { _3571,
                    _544 };
    assign _822 = { _3571,
                    _564 };
    assign _819 = { _3571,
                    _587 };
    assign _795 = { _3571,
                    _532 };
    assign _792 = { _3571,
                    _544 };
    assign _789 = { _3571,
                    _564 };
    assign _786 = { _3571,
                    _539 };
    assign _783 = { _3571,
                    _554 };
    assign _765 = { _3571,
                    _532 };
    assign _545 = { _3571,
                    _544 };
    assign _540 = { _3571,
                    _539 };
    assign _536 = { _3571,
                    _535 };
    assign _541 = _536 + _540;
    assign _546 = _541 + _545;
    assign _548 = _546 < _3574;
    assign _549 = _532 & _548;
    assign _3170 = ~ _549;
    assign _3171 = _532 & _3170;
    assign _3172 = _219 ? _3171 : _532;
    assign _3173 = _529 ? _544 : _3172;
    assign _101 = _3173;
    always @(posedge _207) begin
        if (_221)
            _532 <= _2927;
        else
            _532 <= _101;
    end
    assign _568 = { _3571,
                    _532 };
    assign _591 = { _3571,
                    _544 };
    assign _614 = { _3571,
                    _564 };
    assign _637 = { _3571,
                    _587 };
    assign _660 = { _3571,
                    _610 };
    assign _683 = { _3571,
                    _633 };
    assign _706 = { _3571,
                    _656 };
    assign _729 = { _3571,
                    _679 };
    assign _742 = { _3571,
                    _702 };
    assign _739 = { _3571,
                    _692 };
    assign _737 = { _3571,
                    _715 };
    assign _740 = _737 + _739;
    assign _743 = _740 + _742;
    assign _745 = _743 < _3574;
    assign _746 = _725 & _745;
    assign _3174 = ~ _746;
    assign _3175 = _725 & _3174;
    assign _3176 = _219 ? _3175 : _725;
    assign _3177 = _529 ? _539 : _3176;
    assign _102 = _3177;
    always @(posedge _207) begin
        if (_221)
            _725 <= _2927;
        else
            _725 <= _102;
    end
    assign _726 = { _3571,
                    _725 };
    assign _721 = { _3571,
                    _669 };
    assign _718 = { _3571,
                    _692 };
    assign _716 = { _3571,
                    _715 };
    assign _719 = _716 + _718;
    assign _722 = _719 + _721;
    assign _727 = _722 + _726;
    assign _730 = _727 + _729;
    assign _732 = _730 < _3574;
    assign _733 = _702 & _732;
    assign _3178 = ~ _733;
    assign _3179 = _702 & _3178;
    assign _3180 = _219 ? _3179 : _702;
    assign _3181 = _529 ? _725 : _3180;
    assign _103 = _3181;
    always @(posedge _207) begin
        if (_221)
            _702 <= _2927;
        else
            _702 <= _103;
    end
    assign _703 = { _3571,
                    _702 };
    assign _698 = { _3571,
                    _646 };
    assign _695 = { _3571,
                    _669 };
    assign _693 = { _3571,
                    _692 };
    assign _696 = _693 + _695;
    assign _699 = _696 + _698;
    assign _704 = _699 + _703;
    assign _707 = _704 + _706;
    assign _709 = _707 < _3574;
    assign _710 = _679 & _709;
    assign _3182 = ~ _710;
    assign _3183 = _679 & _3182;
    assign _3184 = _219 ? _3183 : _679;
    assign _3185 = _529 ? _702 : _3184;
    assign _104 = _3185;
    always @(posedge _207) begin
        if (_221)
            _679 <= _2927;
        else
            _679 <= _104;
    end
    assign _680 = { _3571,
                    _679 };
    assign _675 = { _3571,
                    _623 };
    assign _672 = { _3571,
                    _646 };
    assign _670 = { _3571,
                    _669 };
    assign _673 = _670 + _672;
    assign _676 = _673 + _675;
    assign _681 = _676 + _680;
    assign _684 = _681 + _683;
    assign _686 = _684 < _3574;
    assign _687 = _656 & _686;
    assign _3186 = ~ _687;
    assign _3187 = _656 & _3186;
    assign _3188 = _219 ? _3187 : _656;
    assign _3189 = _529 ? _679 : _3188;
    assign _105 = _3189;
    always @(posedge _207) begin
        if (_221)
            _656 <= _2927;
        else
            _656 <= _105;
    end
    assign _657 = { _3571,
                    _656 };
    assign _652 = { _3571,
                    _600 };
    assign _649 = { _3571,
                    _623 };
    assign _647 = { _3571,
                    _646 };
    assign _650 = _647 + _649;
    assign _653 = _650 + _652;
    assign _658 = _653 + _657;
    assign _661 = _658 + _660;
    assign _663 = _661 < _3574;
    assign _664 = _633 & _663;
    assign _3190 = ~ _664;
    assign _3191 = _633 & _3190;
    assign _3192 = _219 ? _3191 : _633;
    assign _3193 = _529 ? _656 : _3192;
    assign _106 = _3193;
    always @(posedge _207) begin
        if (_221)
            _633 <= _2927;
        else
            _633 <= _106;
    end
    assign _634 = { _3571,
                    _633 };
    assign _629 = { _3571,
                    _577 };
    assign _626 = { _3571,
                    _600 };
    assign _624 = { _3571,
                    _623 };
    assign _627 = _624 + _626;
    assign _630 = _627 + _629;
    assign _635 = _630 + _634;
    assign _638 = _635 + _637;
    assign _640 = _638 < _3574;
    assign _641 = _610 & _640;
    assign _3194 = ~ _641;
    assign _3195 = _610 & _3194;
    assign _3196 = _219 ? _3195 : _610;
    assign _3197 = _529 ? _633 : _3196;
    assign _107 = _3197;
    always @(posedge _207) begin
        if (_221)
            _610 <= _2927;
        else
            _610 <= _107;
    end
    assign _611 = { _3571,
                    _610 };
    assign _606 = { _3571,
                    _554 };
    assign _603 = { _3571,
                    _577 };
    assign _601 = { _3571,
                    _600 };
    assign _604 = _601 + _603;
    assign _607 = _604 + _606;
    assign _612 = _607 + _611;
    assign _615 = _612 + _614;
    assign _617 = _615 < _3574;
    assign _618 = _587 & _617;
    assign _3198 = ~ _618;
    assign _3199 = _587 & _3198;
    assign _3200 = _219 ? _3199 : _587;
    assign _3201 = _529 ? _610 : _3200;
    assign _108 = _3201;
    always @(posedge _207) begin
        if (_221)
            _587 <= _2927;
        else
            _587 <= _108;
    end
    assign _588 = { _3571,
                    _587 };
    assign _583 = { _3571,
                    _535 };
    assign _580 = { _3571,
                    _554 };
    assign _578 = { _3571,
                    _577 };
    assign _581 = _578 + _580;
    assign _584 = _581 + _583;
    assign _589 = _584 + _588;
    assign _592 = _589 + _591;
    assign _594 = _592 < _3574;
    assign _595 = _564 & _594;
    assign _3202 = ~ _595;
    assign _3203 = _564 & _3202;
    assign _3204 = _219 ? _3203 : _564;
    assign _3205 = _529 ? _587 : _3204;
    assign _109 = _3205;
    always @(posedge _207) begin
        if (_221)
            _564 <= _2927;
        else
            _564 <= _109;
    end
    assign _565 = { _3571,
                    _564 };
    assign _560 = { _3571,
                    _539 };
    assign _557 = { _3571,
                    _535 };
    assign _555 = { _3571,
                    _554 };
    assign _558 = _555 + _557;
    assign _561 = _558 + _560;
    assign _566 = _561 + _565;
    assign _569 = _566 + _568;
    assign _571 = _569 < _3574;
    assign _572 = _544 & _571;
    assign _3206 = ~ _572;
    assign _3207 = _544 & _3206;
    assign _3208 = _219 ? _3207 : _544;
    assign _3209 = _529 ? _564 : _3208;
    assign _110 = _3209;
    always @(posedge _207) begin
        if (_221)
            _544 <= _2927;
        else
            _544 <= _110;
    end
    assign _762 = { _3571,
                    _544 };
    assign _759 = { _3571,
                    _535 };
    assign _756 = { _3571,
                    _755 };
    assign _752 = { _3571,
                    _751 };
    assign _757 = _752 + _756;
    assign _760 = _757 + _759;
    assign _763 = _760 + _762;
    assign _766 = _763 + _765;
    assign _768 = _766 < _3574;
    assign _769 = _539 & _768;
    assign _3210 = ~ _769;
    assign _3211 = _539 & _3210;
    assign _3212 = _219 ? _3211 : _539;
    assign _3213 = _529 ? _535 : _3212;
    assign _111 = _3213;
    always @(posedge _207) begin
        if (_221)
            _539 <= _2927;
        else
            _539 <= _111;
    end
    assign _1047 = { _3571,
                     _539 };
    assign _1044 = { _3571,
                     _535 };
    assign _1041 = { _3571,
                     _751 };
    assign _1038 = { _3571,
                     _1037 };
    assign _1034 = { _3571,
                     _1033 };
    assign _1039 = _1034 + _1038;
    assign _1042 = _1039 + _1041;
    assign _1045 = _1042 + _1044;
    assign _1048 = _1045 + _1047;
    assign _1050 = _1048 < _3574;
    assign _1051 = _755 & _1050;
    assign _3214 = ~ _1051;
    assign _3215 = _755 & _3214;
    assign _3216 = _219 ? _3215 : _755;
    assign _3217 = _529 ? _751 : _3216;
    assign _112 = _3217;
    always @(posedge _207) begin
        if (_221)
            _755 <= _2927;
        else
            _755 <= _112;
    end
    assign _780 = { _3571,
                    _755 };
    assign _777 = { _3571,
                    _751 };
    assign _775 = { _3571,
                    _774 };
    assign _778 = _775 + _777;
    assign _781 = _778 + _780;
    assign _784 = _781 + _783;
    assign _787 = _784 + _786;
    assign _790 = _787 + _789;
    assign _793 = _790 + _792;
    assign _796 = _793 + _795;
    assign _798 = _796 < _3574;
    assign _799 = _535 & _798;
    assign _3218 = ~ _799;
    assign _3219 = _535 & _3218;
    assign _3220 = _219 ? _3219 : _535;
    assign _3221 = _529 ? _554 : _3220;
    assign _113 = _3221;
    always @(posedge _207) begin
        if (_221)
            _535 <= _2927;
        else
            _535 <= _113;
    end
    assign _816 = { _3571,
                    _535 };
    assign _813 = { _3571,
                    _577 };
    assign _810 = { _3571,
                    _751 };
    assign _807 = { _3571,
                    _774 };
    assign _805 = { _3571,
                    _804 };
    assign _808 = _805 + _807;
    assign _811 = _808 + _810;
    assign _814 = _811 + _813;
    assign _817 = _814 + _816;
    assign _820 = _817 + _819;
    assign _823 = _820 + _822;
    assign _826 = _823 + _825;
    assign _828 = _826 < _3574;
    assign _829 = _554 & _828;
    assign _3222 = ~ _829;
    assign _3223 = _554 & _3222;
    assign _3224 = _219 ? _3223 : _554;
    assign _3225 = _529 ? _577 : _3224;
    assign _114 = _3225;
    always @(posedge _207) begin
        if (_221)
            _554 <= _2927;
        else
            _554 <= _114;
    end
    assign _846 = { _3571,
                    _554 };
    assign _843 = { _3571,
                    _600 };
    assign _840 = { _3571,
                    _774 };
    assign _837 = { _3571,
                    _804 };
    assign _835 = { _3571,
                    _834 };
    assign _838 = _835 + _837;
    assign _841 = _838 + _840;
    assign _844 = _841 + _843;
    assign _847 = _844 + _846;
    assign _850 = _847 + _849;
    assign _853 = _850 + _852;
    assign _856 = _853 + _855;
    assign _858 = _856 < _3574;
    assign _859 = _577 & _858;
    assign _3226 = ~ _859;
    assign _3227 = _577 & _3226;
    assign _3228 = _219 ? _3227 : _577;
    assign _3229 = _529 ? _600 : _3228;
    assign _115 = _3229;
    always @(posedge _207) begin
        if (_221)
            _577 <= _2927;
        else
            _577 <= _115;
    end
    assign _876 = { _3571,
                    _577 };
    assign _873 = { _3571,
                    _623 };
    assign _870 = { _3571,
                    _804 };
    assign _867 = { _3571,
                    _834 };
    assign _865 = { _3571,
                    _864 };
    assign _868 = _865 + _867;
    assign _871 = _868 + _870;
    assign _874 = _871 + _873;
    assign _877 = _874 + _876;
    assign _880 = _877 + _879;
    assign _883 = _880 + _882;
    assign _886 = _883 + _885;
    assign _888 = _886 < _3574;
    assign _889 = _600 & _888;
    assign _3230 = ~ _889;
    assign _3231 = _600 & _3230;
    assign _3232 = _219 ? _3231 : _600;
    assign _3233 = _529 ? _623 : _3232;
    assign _116 = _3233;
    always @(posedge _207) begin
        if (_221)
            _600 <= _2927;
        else
            _600 <= _116;
    end
    assign _906 = { _3571,
                    _600 };
    assign _903 = { _3571,
                    _646 };
    assign _900 = { _3571,
                    _834 };
    assign _897 = { _3571,
                    _864 };
    assign _895 = { _3571,
                    _894 };
    assign _898 = _895 + _897;
    assign _901 = _898 + _900;
    assign _904 = _901 + _903;
    assign _907 = _904 + _906;
    assign _910 = _907 + _909;
    assign _913 = _910 + _912;
    assign _916 = _913 + _915;
    assign _918 = _916 < _3574;
    assign _919 = _623 & _918;
    assign _3234 = ~ _919;
    assign _3235 = _623 & _3234;
    assign _3236 = _219 ? _3235 : _623;
    assign _3237 = _529 ? _646 : _3236;
    assign _117 = _3237;
    always @(posedge _207) begin
        if (_221)
            _623 <= _2927;
        else
            _623 <= _117;
    end
    assign _936 = { _3571,
                    _623 };
    assign _933 = { _3571,
                    _669 };
    assign _930 = { _3571,
                    _864 };
    assign _927 = { _3571,
                    _894 };
    assign _925 = { _3571,
                    _924 };
    assign _928 = _925 + _927;
    assign _931 = _928 + _930;
    assign _934 = _931 + _933;
    assign _937 = _934 + _936;
    assign _940 = _937 + _939;
    assign _943 = _940 + _942;
    assign _946 = _943 + _945;
    assign _948 = _946 < _3574;
    assign _949 = _646 & _948;
    assign _3238 = ~ _949;
    assign _3239 = _646 & _3238;
    assign _3240 = _219 ? _3239 : _646;
    assign _3241 = _529 ? _669 : _3240;
    assign _118 = _3241;
    always @(posedge _207) begin
        if (_221)
            _646 <= _2927;
        else
            _646 <= _118;
    end
    assign _966 = { _3571,
                    _646 };
    assign _963 = { _3571,
                    _692 };
    assign _960 = { _3571,
                    _894 };
    assign _957 = { _3571,
                    _924 };
    assign _955 = { _3571,
                    _954 };
    assign _958 = _955 + _957;
    assign _961 = _958 + _960;
    assign _964 = _961 + _963;
    assign _967 = _964 + _966;
    assign _970 = _967 + _969;
    assign _973 = _970 + _972;
    assign _976 = _973 + _975;
    assign _978 = _976 < _3574;
    assign _979 = _669 & _978;
    assign _3242 = ~ _979;
    assign _3243 = _669 & _3242;
    assign _3244 = _219 ? _3243 : _669;
    assign _3245 = _529 ? _692 : _3244;
    assign _119 = _3245;
    always @(posedge _207) begin
        if (_221)
            _669 <= _2927;
        else
            _669 <= _119;
    end
    assign _996 = { _3571,
                    _669 };
    assign _993 = { _3571,
                    _715 };
    assign _990 = { _3571,
                    _924 };
    assign _987 = { _3571,
                    _954 };
    assign _985 = { _3571,
                    _984 };
    assign _988 = _985 + _987;
    assign _991 = _988 + _990;
    assign _994 = _991 + _993;
    assign _997 = _994 + _996;
    assign _1000 = _997 + _999;
    assign _1003 = _1000 + _1002;
    assign _1006 = _1003 + _1005;
    assign _1008 = _1006 < _3574;
    assign _1009 = _692 & _1008;
    assign _3246 = ~ _1009;
    assign _3247 = _692 & _3246;
    assign _3248 = _219 ? _3247 : _692;
    assign _3249 = _529 ? _715 : _3248;
    assign _120 = _3249;
    always @(posedge _207) begin
        if (_221)
            _692 <= _2927;
        else
            _692 <= _120;
    end
    assign _1018 = { _3571,
                     _692 };
    assign _1015 = { _3571,
                     _954 };
    assign _1013 = { _3571,
                     _984 };
    assign _1016 = _1013 + _1015;
    assign _1019 = _1016 + _1018;
    assign _1022 = _1019 + _1021;
    assign _1025 = _1022 + _1024;
    assign _1027 = _1025 < _3574;
    assign _1028 = _715 & _1027;
    assign _3250 = ~ _1028;
    assign _3251 = _715 & _3250;
    assign _3252 = _219 ? _3251 : _715;
    assign _3253 = _529 ? _755 : _3252;
    assign _121 = _3253;
    always @(posedge _207) begin
        if (_221)
            _715 <= _2927;
        else
            _715 <= _121;
    end
    assign _1303 = { _3571,
                     _715 };
    assign _1300 = { _3571,
                     _954 };
    assign _1297 = { _3571,
                     _1236 };
    assign _1295 = { _3571,
                     _1266 };
    assign _1298 = _1295 + _1297;
    assign _1301 = _1298 + _1300;
    assign _1304 = _1301 + _1303;
    assign _1307 = _1304 + _1306;
    assign _1309 = _1307 < _3574;
    assign _1310 = _984 & _1309;
    assign _3254 = ~ _1310;
    assign _3255 = _984 & _3254;
    assign _3256 = _219 ? _3255 : _984;
    assign _3257 = _529 ? _1037 : _3256;
    assign _122 = _3257;
    always @(posedge _207) begin
        if (_221)
            _984 <= _2927;
        else
            _984 <= _122;
    end
    assign _1275 = { _3571,
                     _984 };
    assign _1272 = { _3571,
                     _1206 };
    assign _1269 = { _3571,
                     _1236 };
    assign _1267 = { _3571,
                     _1266 };
    assign _1270 = _1267 + _1269;
    assign _1273 = _1270 + _1272;
    assign _1276 = _1273 + _1275;
    assign _1279 = _1276 + _1278;
    assign _1282 = _1279 + _1281;
    assign _1285 = _1282 + _1284;
    assign _1288 = _1285 + _1287;
    assign _1290 = _1288 < _3574;
    assign _1291 = _954 & _1290;
    assign _3258 = ~ _1291;
    assign _3259 = _954 & _3258;
    assign _3260 = _219 ? _3259 : _954;
    assign _3261 = _529 ? _984 : _3260;
    assign _123 = _3261;
    always @(posedge _207) begin
        if (_221)
            _954 <= _2927;
        else
            _954 <= _123;
    end
    assign _1245 = { _3571,
                     _954 };
    assign _1242 = { _3571,
                     _1176 };
    assign _1239 = { _3571,
                     _1206 };
    assign _1237 = { _3571,
                     _1236 };
    assign _1240 = _1237 + _1239;
    assign _1243 = _1240 + _1242;
    assign _1246 = _1243 + _1245;
    assign _1249 = _1246 + _1248;
    assign _1252 = _1249 + _1251;
    assign _1255 = _1252 + _1254;
    assign _1258 = _1255 + _1257;
    assign _1260 = _1258 < _3574;
    assign _1261 = _924 & _1260;
    assign _3262 = ~ _1261;
    assign _3263 = _924 & _3262;
    assign _3264 = _219 ? _3263 : _924;
    assign _3265 = _529 ? _954 : _3264;
    assign _124 = _3265;
    always @(posedge _207) begin
        if (_221)
            _924 <= _2927;
        else
            _924 <= _124;
    end
    assign _1215 = { _3571,
                     _924 };
    assign _1212 = { _3571,
                     _1146 };
    assign _1209 = { _3571,
                     _1176 };
    assign _1207 = { _3571,
                     _1206 };
    assign _1210 = _1207 + _1209;
    assign _1213 = _1210 + _1212;
    assign _1216 = _1213 + _1215;
    assign _1219 = _1216 + _1218;
    assign _1222 = _1219 + _1221;
    assign _1225 = _1222 + _1224;
    assign _1228 = _1225 + _1227;
    assign _1230 = _1228 < _3574;
    assign _1231 = _894 & _1230;
    assign _3266 = ~ _1231;
    assign _3267 = _894 & _3266;
    assign _3268 = _219 ? _3267 : _894;
    assign _3269 = _529 ? _924 : _3268;
    assign _125 = _3269;
    always @(posedge _207) begin
        if (_221)
            _894 <= _2927;
        else
            _894 <= _125;
    end
    assign _1185 = { _3571,
                     _894 };
    assign _1182 = { _3571,
                     _1116 };
    assign _1179 = { _3571,
                     _1146 };
    assign _1177 = { _3571,
                     _1176 };
    assign _1180 = _1177 + _1179;
    assign _1183 = _1180 + _1182;
    assign _1186 = _1183 + _1185;
    assign _1189 = _1186 + _1188;
    assign _1192 = _1189 + _1191;
    assign _1195 = _1192 + _1194;
    assign _1198 = _1195 + _1197;
    assign _1200 = _1198 < _3574;
    assign _1201 = _864 & _1200;
    assign _3270 = ~ _1201;
    assign _3271 = _864 & _3270;
    assign _3272 = _219 ? _3271 : _864;
    assign _3273 = _529 ? _894 : _3272;
    assign _126 = _3273;
    always @(posedge _207) begin
        if (_221)
            _864 <= _2927;
        else
            _864 <= _126;
    end
    assign _1155 = { _3571,
                     _864 };
    assign _1152 = { _3571,
                     _1086 };
    assign _1149 = { _3571,
                     _1116 };
    assign _1147 = { _3571,
                     _1146 };
    assign _1150 = _1147 + _1149;
    assign _1153 = _1150 + _1152;
    assign _1156 = _1153 + _1155;
    assign _1159 = _1156 + _1158;
    assign _1162 = _1159 + _1161;
    assign _1165 = _1162 + _1164;
    assign _1168 = _1165 + _1167;
    assign _1170 = _1168 < _3574;
    assign _1171 = _834 & _1170;
    assign _3274 = ~ _1171;
    assign _3275 = _834 & _3274;
    assign _3276 = _219 ? _3275 : _834;
    assign _3277 = _529 ? _864 : _3276;
    assign _127 = _3277;
    always @(posedge _207) begin
        if (_221)
            _834 <= _2927;
        else
            _834 <= _127;
    end
    assign _1125 = { _3571,
                     _834 };
    assign _1122 = { _3571,
                     _1056 };
    assign _1119 = { _3571,
                     _1086 };
    assign _1117 = { _3571,
                     _1116 };
    assign _1120 = _1117 + _1119;
    assign _1123 = _1120 + _1122;
    assign _1126 = _1123 + _1125;
    assign _1129 = _1126 + _1128;
    assign _1132 = _1129 + _1131;
    assign _1135 = _1132 + _1134;
    assign _1138 = _1135 + _1137;
    assign _1140 = _1138 < _3574;
    assign _1141 = _804 & _1140;
    assign _3278 = ~ _1141;
    assign _3279 = _804 & _3278;
    assign _3280 = _219 ? _3279 : _804;
    assign _3281 = _529 ? _834 : _3280;
    assign _128 = _3281;
    always @(posedge _207) begin
        if (_221)
            _804 <= _2927;
        else
            _804 <= _128;
    end
    assign _1095 = { _3571,
                     _804 };
    assign _1092 = { _3571,
                     _1033 };
    assign _1089 = { _3571,
                     _1056 };
    assign _1087 = { _3571,
                     _1086 };
    assign _1090 = _1087 + _1089;
    assign _1093 = _1090 + _1092;
    assign _1096 = _1093 + _1095;
    assign _1099 = _1096 + _1098;
    assign _1102 = _1099 + _1101;
    assign _1105 = _1102 + _1104;
    assign _1108 = _1105 + _1107;
    assign _1110 = _1108 < _3574;
    assign _1111 = _774 & _1110;
    assign _3282 = ~ _1111;
    assign _3283 = _774 & _3282;
    assign _3284 = _219 ? _3283 : _774;
    assign _3285 = _529 ? _804 : _3284;
    assign _129 = _3285;
    always @(posedge _207) begin
        if (_221)
            _774 <= _2927;
        else
            _774 <= _129;
    end
    assign _1065 = { _3571,
                     _774 };
    assign _1062 = { _3571,
                     _1037 };
    assign _1059 = { _3571,
                     _1033 };
    assign _1057 = { _3571,
                     _1056 };
    assign _1060 = _1057 + _1059;
    assign _1063 = _1060 + _1062;
    assign _1066 = _1063 + _1065;
    assign _1069 = _1066 + _1068;
    assign _1072 = _1069 + _1071;
    assign _1075 = _1072 + _1074;
    assign _1078 = _1075 + _1077;
    assign _1080 = _1078 < _3574;
    assign _1081 = _751 & _1080;
    assign _3286 = ~ _1081;
    assign _3287 = _751 & _3286;
    assign _3288 = _219 ? _3287 : _751;
    assign _3289 = _529 ? _774 : _3288;
    assign _130 = _3289;
    always @(posedge _207) begin
        if (_221)
            _751 <= _2927;
        else
            _751 <= _130;
    end
    assign _1326 = { _3571,
                     _751 };
    assign _1323 = { _3571,
                     _1033 };
    assign _1320 = { _3571,
                     _1319 };
    assign _1316 = { _3571,
                     _1315 };
    assign _1321 = _1316 + _1320;
    assign _1324 = _1321 + _1323;
    assign _1327 = _1324 + _1326;
    assign _1330 = _1327 + _1329;
    assign _1332 = _1330 < _3574;
    assign _1333 = _1037 & _1332;
    assign _3290 = ~ _1333;
    assign _3291 = _1037 & _3290;
    assign _3292 = _219 ? _3291 : _1037;
    assign _3293 = _529 ? _1033 : _3292;
    assign _131 = _3293;
    always @(posedge _207) begin
        if (_221)
            _1037 <= _2927;
        else
            _1037 <= _131;
    end
    assign _1611 = { _3571,
                     _1037 };
    assign _1608 = { _3571,
                     _1033 };
    assign _1605 = { _3571,
                     _1315 };
    assign _1602 = { _3571,
                     _1601 };
    assign _1598 = { _3571,
                     _1597 };
    assign _1603 = _1598 + _1602;
    assign _1606 = _1603 + _1605;
    assign _1609 = _1606 + _1608;
    assign _1612 = _1609 + _1611;
    assign _1614 = _1612 < _3574;
    assign _1615 = _1319 & _1614;
    assign _3294 = ~ _1615;
    assign _3295 = _1319 & _3294;
    assign _3296 = _219 ? _3295 : _1319;
    assign _3297 = _529 ? _1315 : _3296;
    assign _132 = _3297;
    always @(posedge _207) begin
        if (_221)
            _1319 <= _2927;
        else
            _1319 <= _132;
    end
    assign _1344 = { _3571,
                     _1319 };
    assign _1341 = { _3571,
                     _1315 };
    assign _1339 = { _3571,
                     _1338 };
    assign _1342 = _1339 + _1341;
    assign _1345 = _1342 + _1344;
    assign _1348 = _1345 + _1347;
    assign _1351 = _1348 + _1350;
    assign _1354 = _1351 + _1353;
    assign _1357 = _1354 + _1356;
    assign _1360 = _1357 + _1359;
    assign _1362 = _1360 < _3574;
    assign _1363 = _1033 & _1362;
    assign _3298 = ~ _1363;
    assign _3299 = _1033 & _3298;
    assign _3300 = _219 ? _3299 : _1033;
    assign _3301 = _529 ? _1056 : _3300;
    assign _133 = _3301;
    always @(posedge _207) begin
        if (_221)
            _1033 <= _2927;
        else
            _1033 <= _133;
    end
    assign _1380 = { _3571,
                     _1033 };
    assign _1377 = { _3571,
                     _1086 };
    assign _1374 = { _3571,
                     _1315 };
    assign _1371 = { _3571,
                     _1338 };
    assign _1369 = { _3571,
                     _1368 };
    assign _1372 = _1369 + _1371;
    assign _1375 = _1372 + _1374;
    assign _1378 = _1375 + _1377;
    assign _1381 = _1378 + _1380;
    assign _1384 = _1381 + _1383;
    assign _1387 = _1384 + _1386;
    assign _1390 = _1387 + _1389;
    assign _1392 = _1390 < _3574;
    assign _1393 = _1056 & _1392;
    assign _3302 = ~ _1393;
    assign _3303 = _1056 & _3302;
    assign _3304 = _219 ? _3303 : _1056;
    assign _3305 = _529 ? _1086 : _3304;
    assign _134 = _3305;
    always @(posedge _207) begin
        if (_221)
            _1056 <= _2927;
        else
            _1056 <= _134;
    end
    assign _1410 = { _3571,
                     _1056 };
    assign _1407 = { _3571,
                     _1116 };
    assign _1404 = { _3571,
                     _1338 };
    assign _1401 = { _3571,
                     _1368 };
    assign _1399 = { _3571,
                     _1398 };
    assign _1402 = _1399 + _1401;
    assign _1405 = _1402 + _1404;
    assign _1408 = _1405 + _1407;
    assign _1411 = _1408 + _1410;
    assign _1414 = _1411 + _1413;
    assign _1417 = _1414 + _1416;
    assign _1420 = _1417 + _1419;
    assign _1422 = _1420 < _3574;
    assign _1423 = _1086 & _1422;
    assign _3306 = ~ _1423;
    assign _3307 = _1086 & _3306;
    assign _3308 = _219 ? _3307 : _1086;
    assign _3309 = _529 ? _1116 : _3308;
    assign _135 = _3309;
    always @(posedge _207) begin
        if (_221)
            _1086 <= _2927;
        else
            _1086 <= _135;
    end
    assign _1440 = { _3571,
                     _1086 };
    assign _1437 = { _3571,
                     _1146 };
    assign _1434 = { _3571,
                     _1368 };
    assign _1431 = { _3571,
                     _1398 };
    assign _1429 = { _3571,
                     _1428 };
    assign _1432 = _1429 + _1431;
    assign _1435 = _1432 + _1434;
    assign _1438 = _1435 + _1437;
    assign _1441 = _1438 + _1440;
    assign _1444 = _1441 + _1443;
    assign _1447 = _1444 + _1446;
    assign _1450 = _1447 + _1449;
    assign _1452 = _1450 < _3574;
    assign _1453 = _1116 & _1452;
    assign _3310 = ~ _1453;
    assign _3311 = _1116 & _3310;
    assign _3312 = _219 ? _3311 : _1116;
    assign _3313 = _529 ? _1146 : _3312;
    assign _136 = _3313;
    always @(posedge _207) begin
        if (_221)
            _1116 <= _2927;
        else
            _1116 <= _136;
    end
    assign _1470 = { _3571,
                     _1116 };
    assign _1467 = { _3571,
                     _1176 };
    assign _1464 = { _3571,
                     _1398 };
    assign _1461 = { _3571,
                     _1428 };
    assign _1459 = { _3571,
                     _1458 };
    assign _1462 = _1459 + _1461;
    assign _1465 = _1462 + _1464;
    assign _1468 = _1465 + _1467;
    assign _1471 = _1468 + _1470;
    assign _1474 = _1471 + _1473;
    assign _1477 = _1474 + _1476;
    assign _1480 = _1477 + _1479;
    assign _1482 = _1480 < _3574;
    assign _1483 = _1146 & _1482;
    assign _3314 = ~ _1483;
    assign _3315 = _1146 & _3314;
    assign _3316 = _219 ? _3315 : _1146;
    assign _3317 = _529 ? _1176 : _3316;
    assign _137 = _3317;
    always @(posedge _207) begin
        if (_221)
            _1146 <= _2927;
        else
            _1146 <= _137;
    end
    assign _1500 = { _3571,
                     _1146 };
    assign _1497 = { _3571,
                     _1206 };
    assign _1494 = { _3571,
                     _1428 };
    assign _1491 = { _3571,
                     _1458 };
    assign _1489 = { _3571,
                     _1488 };
    assign _1492 = _1489 + _1491;
    assign _1495 = _1492 + _1494;
    assign _1498 = _1495 + _1497;
    assign _1501 = _1498 + _1500;
    assign _1504 = _1501 + _1503;
    assign _1507 = _1504 + _1506;
    assign _1510 = _1507 + _1509;
    assign _1512 = _1510 < _3574;
    assign _1513 = _1176 & _1512;
    assign _3318 = ~ _1513;
    assign _3319 = _1176 & _3318;
    assign _3320 = _219 ? _3319 : _1176;
    assign _3321 = _529 ? _1206 : _3320;
    assign _138 = _3321;
    always @(posedge _207) begin
        if (_221)
            _1176 <= _2927;
        else
            _1176 <= _138;
    end
    assign _1530 = { _3571,
                     _1176 };
    assign _1527 = { _3571,
                     _1236 };
    assign _1524 = { _3571,
                     _1458 };
    assign _1521 = { _3571,
                     _1488 };
    assign _1519 = { _3571,
                     _1518 };
    assign _1522 = _1519 + _1521;
    assign _1525 = _1522 + _1524;
    assign _1528 = _1525 + _1527;
    assign _1531 = _1528 + _1530;
    assign _1534 = _1531 + _1533;
    assign _1537 = _1534 + _1536;
    assign _1540 = _1537 + _1539;
    assign _1542 = _1540 < _3574;
    assign _1543 = _1206 & _1542;
    assign _3322 = ~ _1543;
    assign _3323 = _1206 & _3322;
    assign _3324 = _219 ? _3323 : _1206;
    assign _3325 = _529 ? _1236 : _3324;
    assign _139 = _3325;
    always @(posedge _207) begin
        if (_221)
            _1206 <= _2927;
        else
            _1206 <= _139;
    end
    assign _1560 = { _3571,
                     _1206 };
    assign _1557 = { _3571,
                     _1266 };
    assign _1554 = { _3571,
                     _1488 };
    assign _1551 = { _3571,
                     _1518 };
    assign _1549 = { _3571,
                     _1548 };
    assign _1552 = _1549 + _1551;
    assign _1555 = _1552 + _1554;
    assign _1558 = _1555 + _1557;
    assign _1561 = _1558 + _1560;
    assign _1564 = _1561 + _1563;
    assign _1567 = _1564 + _1566;
    assign _1570 = _1567 + _1569;
    assign _1572 = _1570 < _3574;
    assign _1573 = _1236 & _1572;
    assign _3326 = ~ _1573;
    assign _3327 = _1236 & _3326;
    assign _3328 = _219 ? _3327 : _1236;
    assign _3329 = _529 ? _1266 : _3328;
    assign _140 = _3329;
    always @(posedge _207) begin
        if (_221)
            _1236 <= _2927;
        else
            _1236 <= _140;
    end
    assign _1582 = { _3571,
                     _1236 };
    assign _1579 = { _3571,
                     _1518 };
    assign _1577 = { _3571,
                     _1548 };
    assign _1580 = _1577 + _1579;
    assign _1583 = _1580 + _1582;
    assign _1586 = _1583 + _1585;
    assign _1589 = _1586 + _1588;
    assign _1591 = _1589 < _3574;
    assign _1592 = _1266 & _1591;
    assign _3330 = ~ _1592;
    assign _3331 = _1266 & _3330;
    assign _3332 = _219 ? _3331 : _1266;
    assign _3333 = _529 ? _1319 : _3332;
    assign _141 = _3333;
    always @(posedge _207) begin
        if (_221)
            _1266 <= _2927;
        else
            _1266 <= _141;
    end
    assign _1867 = { _3571,
                     _1266 };
    assign _1864 = { _3571,
                     _1518 };
    assign _1861 = { _3571,
                     _1800 };
    assign _1859 = { _3571,
                     _1830 };
    assign _1862 = _1859 + _1861;
    assign _1865 = _1862 + _1864;
    assign _1868 = _1865 + _1867;
    assign _1871 = _1868 + _1870;
    assign _1873 = _1871 < _3574;
    assign _1874 = _1548 & _1873;
    assign _3334 = ~ _1874;
    assign _3335 = _1548 & _3334;
    assign _3336 = _219 ? _3335 : _1548;
    assign _3337 = _529 ? _1601 : _3336;
    assign _142 = _3337;
    always @(posedge _207) begin
        if (_221)
            _1548 <= _2927;
        else
            _1548 <= _142;
    end
    assign _1839 = { _3571,
                     _1548 };
    assign _1836 = { _3571,
                     _1770 };
    assign _1833 = { _3571,
                     _1800 };
    assign _1831 = { _3571,
                     _1830 };
    assign _1834 = _1831 + _1833;
    assign _1837 = _1834 + _1836;
    assign _1840 = _1837 + _1839;
    assign _1843 = _1840 + _1842;
    assign _1846 = _1843 + _1845;
    assign _1849 = _1846 + _1848;
    assign _1852 = _1849 + _1851;
    assign _1854 = _1852 < _3574;
    assign _1855 = _1518 & _1854;
    assign _3338 = ~ _1855;
    assign _3339 = _1518 & _3338;
    assign _3340 = _219 ? _3339 : _1518;
    assign _3341 = _529 ? _1548 : _3340;
    assign _143 = _3341;
    always @(posedge _207) begin
        if (_221)
            _1518 <= _2927;
        else
            _1518 <= _143;
    end
    assign _1809 = { _3571,
                     _1518 };
    assign _1806 = { _3571,
                     _1740 };
    assign _1803 = { _3571,
                     _1770 };
    assign _1801 = { _3571,
                     _1800 };
    assign _1804 = _1801 + _1803;
    assign _1807 = _1804 + _1806;
    assign _1810 = _1807 + _1809;
    assign _1813 = _1810 + _1812;
    assign _1816 = _1813 + _1815;
    assign _1819 = _1816 + _1818;
    assign _1822 = _1819 + _1821;
    assign _1824 = _1822 < _3574;
    assign _1825 = _1488 & _1824;
    assign _3342 = ~ _1825;
    assign _3343 = _1488 & _3342;
    assign _3344 = _219 ? _3343 : _1488;
    assign _3345 = _529 ? _1518 : _3344;
    assign _144 = _3345;
    always @(posedge _207) begin
        if (_221)
            _1488 <= _2927;
        else
            _1488 <= _144;
    end
    assign _1779 = { _3571,
                     _1488 };
    assign _1776 = { _3571,
                     _1710 };
    assign _1773 = { _3571,
                     _1740 };
    assign _1771 = { _3571,
                     _1770 };
    assign _1774 = _1771 + _1773;
    assign _1777 = _1774 + _1776;
    assign _1780 = _1777 + _1779;
    assign _1783 = _1780 + _1782;
    assign _1786 = _1783 + _1785;
    assign _1789 = _1786 + _1788;
    assign _1792 = _1789 + _1791;
    assign _1794 = _1792 < _3574;
    assign _1795 = _1458 & _1794;
    assign _3346 = ~ _1795;
    assign _3347 = _1458 & _3346;
    assign _3348 = _219 ? _3347 : _1458;
    assign _3349 = _529 ? _1488 : _3348;
    assign _145 = _3349;
    always @(posedge _207) begin
        if (_221)
            _1458 <= _2927;
        else
            _1458 <= _145;
    end
    assign _1749 = { _3571,
                     _1458 };
    assign _1746 = { _3571,
                     _1680 };
    assign _1743 = { _3571,
                     _1710 };
    assign _1741 = { _3571,
                     _1740 };
    assign _1744 = _1741 + _1743;
    assign _1747 = _1744 + _1746;
    assign _1750 = _1747 + _1749;
    assign _1753 = _1750 + _1752;
    assign _1756 = _1753 + _1755;
    assign _1759 = _1756 + _1758;
    assign _1762 = _1759 + _1761;
    assign _1764 = _1762 < _3574;
    assign _1765 = _1428 & _1764;
    assign _3350 = ~ _1765;
    assign _3351 = _1428 & _3350;
    assign _3352 = _219 ? _3351 : _1428;
    assign _3353 = _529 ? _1458 : _3352;
    assign _146 = _3353;
    always @(posedge _207) begin
        if (_221)
            _1428 <= _2927;
        else
            _1428 <= _146;
    end
    assign _1719 = { _3571,
                     _1428 };
    assign _1716 = { _3571,
                     _1650 };
    assign _1713 = { _3571,
                     _1680 };
    assign _1711 = { _3571,
                     _1710 };
    assign _1714 = _1711 + _1713;
    assign _1717 = _1714 + _1716;
    assign _1720 = _1717 + _1719;
    assign _1723 = _1720 + _1722;
    assign _1726 = _1723 + _1725;
    assign _1729 = _1726 + _1728;
    assign _1732 = _1729 + _1731;
    assign _1734 = _1732 < _3574;
    assign _1735 = _1398 & _1734;
    assign _3354 = ~ _1735;
    assign _3355 = _1398 & _3354;
    assign _3356 = _219 ? _3355 : _1398;
    assign _3357 = _529 ? _1428 : _3356;
    assign _147 = _3357;
    always @(posedge _207) begin
        if (_221)
            _1398 <= _2927;
        else
            _1398 <= _147;
    end
    assign _1689 = { _3571,
                     _1398 };
    assign _1686 = { _3571,
                     _1620 };
    assign _1683 = { _3571,
                     _1650 };
    assign _1681 = { _3571,
                     _1680 };
    assign _1684 = _1681 + _1683;
    assign _1687 = _1684 + _1686;
    assign _1690 = _1687 + _1689;
    assign _1693 = _1690 + _1692;
    assign _1696 = _1693 + _1695;
    assign _1699 = _1696 + _1698;
    assign _1702 = _1699 + _1701;
    assign _1704 = _1702 < _3574;
    assign _1705 = _1368 & _1704;
    assign _3358 = ~ _1705;
    assign _3359 = _1368 & _3358;
    assign _3360 = _219 ? _3359 : _1368;
    assign _3361 = _529 ? _1398 : _3360;
    assign _148 = _3361;
    always @(posedge _207) begin
        if (_221)
            _1368 <= _2927;
        else
            _1368 <= _148;
    end
    assign _1659 = { _3571,
                     _1368 };
    assign _1656 = { _3571,
                     _1597 };
    assign _1653 = { _3571,
                     _1620 };
    assign _1651 = { _3571,
                     _1650 };
    assign _1654 = _1651 + _1653;
    assign _1657 = _1654 + _1656;
    assign _1660 = _1657 + _1659;
    assign _1663 = _1660 + _1662;
    assign _1666 = _1663 + _1665;
    assign _1669 = _1666 + _1668;
    assign _1672 = _1669 + _1671;
    assign _1674 = _1672 < _3574;
    assign _1675 = _1338 & _1674;
    assign _3362 = ~ _1675;
    assign _3363 = _1338 & _3362;
    assign _3364 = _219 ? _3363 : _1338;
    assign _3365 = _529 ? _1368 : _3364;
    assign _149 = _3365;
    always @(posedge _207) begin
        if (_221)
            _1338 <= _2927;
        else
            _1338 <= _149;
    end
    assign _1629 = { _3571,
                     _1338 };
    assign _1626 = { _3571,
                     _1601 };
    assign _1623 = { _3571,
                     _1597 };
    assign _1621 = { _3571,
                     _1620 };
    assign _1624 = _1621 + _1623;
    assign _1627 = _1624 + _1626;
    assign _1630 = _1627 + _1629;
    assign _1633 = _1630 + _1632;
    assign _1636 = _1633 + _1635;
    assign _1639 = _1636 + _1638;
    assign _1642 = _1639 + _1641;
    assign _1644 = _1642 < _3574;
    assign _1645 = _1315 & _1644;
    assign _3366 = ~ _1645;
    assign _3367 = _1315 & _3366;
    assign _3368 = _219 ? _3367 : _1315;
    assign _3369 = _529 ? _1338 : _3368;
    assign _150 = _3369;
    always @(posedge _207) begin
        if (_221)
            _1315 <= _2927;
        else
            _1315 <= _150;
    end
    assign _1890 = { _3571,
                     _1315 };
    assign _1887 = { _3571,
                     _1597 };
    assign _1884 = { _3571,
                     _1883 };
    assign _1880 = { _3571,
                     _1879 };
    assign _1885 = _1880 + _1884;
    assign _1888 = _1885 + _1887;
    assign _1891 = _1888 + _1890;
    assign _1894 = _1891 + _1893;
    assign _1896 = _1894 < _3574;
    assign _1897 = _1601 & _1896;
    assign _3370 = ~ _1897;
    assign _3371 = _1601 & _3370;
    assign _3372 = _219 ? _3371 : _1601;
    assign _3373 = _529 ? _1597 : _3372;
    assign _151 = _3373;
    always @(posedge _207) begin
        if (_221)
            _1601 <= _2927;
        else
            _1601 <= _151;
    end
    assign _2175 = { _3571,
                     _1601 };
    assign _2172 = { _3571,
                     _1597 };
    assign _2169 = { _3571,
                     _1879 };
    assign _2166 = { _3571,
                     _2165 };
    assign _2162 = { _3571,
                     _2161 };
    assign _2167 = _2162 + _2166;
    assign _2170 = _2167 + _2169;
    assign _2173 = _2170 + _2172;
    assign _2176 = _2173 + _2175;
    assign _2178 = _2176 < _3574;
    assign _2179 = _1883 & _2178;
    assign _3374 = ~ _2179;
    assign _3375 = _1883 & _3374;
    assign _3376 = _219 ? _3375 : _1883;
    assign _3377 = _529 ? _1879 : _3376;
    assign _152 = _3377;
    always @(posedge _207) begin
        if (_221)
            _1883 <= _2927;
        else
            _1883 <= _152;
    end
    assign _1908 = { _3571,
                     _1883 };
    assign _1905 = { _3571,
                     _1879 };
    assign _1903 = { _3571,
                     _1902 };
    assign _1906 = _1903 + _1905;
    assign _1909 = _1906 + _1908;
    assign _1912 = _1909 + _1911;
    assign _1915 = _1912 + _1914;
    assign _1918 = _1915 + _1917;
    assign _1921 = _1918 + _1920;
    assign _1924 = _1921 + _1923;
    assign _1926 = _1924 < _3574;
    assign _1927 = _1597 & _1926;
    assign _3378 = ~ _1927;
    assign _3379 = _1597 & _3378;
    assign _3380 = _219 ? _3379 : _1597;
    assign _3381 = _529 ? _1620 : _3380;
    assign _153 = _3381;
    always @(posedge _207) begin
        if (_221)
            _1597 <= _2927;
        else
            _1597 <= _153;
    end
    assign _1944 = { _3571,
                     _1597 };
    assign _1941 = { _3571,
                     _1650 };
    assign _1938 = { _3571,
                     _1879 };
    assign _1935 = { _3571,
                     _1902 };
    assign _1933 = { _3571,
                     _1932 };
    assign _1936 = _1933 + _1935;
    assign _1939 = _1936 + _1938;
    assign _1942 = _1939 + _1941;
    assign _1945 = _1942 + _1944;
    assign _1948 = _1945 + _1947;
    assign _1951 = _1948 + _1950;
    assign _1954 = _1951 + _1953;
    assign _1956 = _1954 < _3574;
    assign _1957 = _1620 & _1956;
    assign _3382 = ~ _1957;
    assign _3383 = _1620 & _3382;
    assign _3384 = _219 ? _3383 : _1620;
    assign _3385 = _529 ? _1650 : _3384;
    assign _154 = _3385;
    always @(posedge _207) begin
        if (_221)
            _1620 <= _2927;
        else
            _1620 <= _154;
    end
    assign _1974 = { _3571,
                     _1620 };
    assign _1971 = { _3571,
                     _1680 };
    assign _1968 = { _3571,
                     _1902 };
    assign _1965 = { _3571,
                     _1932 };
    assign _1963 = { _3571,
                     _1962 };
    assign _1966 = _1963 + _1965;
    assign _1969 = _1966 + _1968;
    assign _1972 = _1969 + _1971;
    assign _1975 = _1972 + _1974;
    assign _1978 = _1975 + _1977;
    assign _1981 = _1978 + _1980;
    assign _1984 = _1981 + _1983;
    assign _1986 = _1984 < _3574;
    assign _1987 = _1650 & _1986;
    assign _3386 = ~ _1987;
    assign _3387 = _1650 & _3386;
    assign _3388 = _219 ? _3387 : _1650;
    assign _3389 = _529 ? _1680 : _3388;
    assign _155 = _3389;
    always @(posedge _207) begin
        if (_221)
            _1650 <= _2927;
        else
            _1650 <= _155;
    end
    assign _2004 = { _3571,
                     _1650 };
    assign _2001 = { _3571,
                     _1710 };
    assign _1998 = { _3571,
                     _1932 };
    assign _1995 = { _3571,
                     _1962 };
    assign _1993 = { _3571,
                     _1992 };
    assign _1996 = _1993 + _1995;
    assign _1999 = _1996 + _1998;
    assign _2002 = _1999 + _2001;
    assign _2005 = _2002 + _2004;
    assign _2008 = _2005 + _2007;
    assign _2011 = _2008 + _2010;
    assign _2014 = _2011 + _2013;
    assign _2016 = _2014 < _3574;
    assign _2017 = _1680 & _2016;
    assign _3390 = ~ _2017;
    assign _3391 = _1680 & _3390;
    assign _3392 = _219 ? _3391 : _1680;
    assign _3393 = _529 ? _1710 : _3392;
    assign _156 = _3393;
    always @(posedge _207) begin
        if (_221)
            _1680 <= _2927;
        else
            _1680 <= _156;
    end
    assign _2034 = { _3571,
                     _1680 };
    assign _2031 = { _3571,
                     _1740 };
    assign _2028 = { _3571,
                     _1962 };
    assign _2025 = { _3571,
                     _1992 };
    assign _2023 = { _3571,
                     _2022 };
    assign _2026 = _2023 + _2025;
    assign _2029 = _2026 + _2028;
    assign _2032 = _2029 + _2031;
    assign _2035 = _2032 + _2034;
    assign _2038 = _2035 + _2037;
    assign _2041 = _2038 + _2040;
    assign _2044 = _2041 + _2043;
    assign _2046 = _2044 < _3574;
    assign _2047 = _1710 & _2046;
    assign _3394 = ~ _2047;
    assign _3395 = _1710 & _3394;
    assign _3396 = _219 ? _3395 : _1710;
    assign _3397 = _529 ? _1740 : _3396;
    assign _157 = _3397;
    always @(posedge _207) begin
        if (_221)
            _1710 <= _2927;
        else
            _1710 <= _157;
    end
    assign _2064 = { _3571,
                     _1710 };
    assign _2061 = { _3571,
                     _1770 };
    assign _2058 = { _3571,
                     _1992 };
    assign _2055 = { _3571,
                     _2022 };
    assign _2053 = { _3571,
                     _2052 };
    assign _2056 = _2053 + _2055;
    assign _2059 = _2056 + _2058;
    assign _2062 = _2059 + _2061;
    assign _2065 = _2062 + _2064;
    assign _2068 = _2065 + _2067;
    assign _2071 = _2068 + _2070;
    assign _2074 = _2071 + _2073;
    assign _2076 = _2074 < _3574;
    assign _2077 = _1740 & _2076;
    assign _3398 = ~ _2077;
    assign _3399 = _1740 & _3398;
    assign _3400 = _219 ? _3399 : _1740;
    assign _3401 = _529 ? _1770 : _3400;
    assign _158 = _3401;
    always @(posedge _207) begin
        if (_221)
            _1740 <= _2927;
        else
            _1740 <= _158;
    end
    assign _2094 = { _3571,
                     _1740 };
    assign _2091 = { _3571,
                     _1800 };
    assign _2088 = { _3571,
                     _2022 };
    assign _2085 = { _3571,
                     _2052 };
    assign _2083 = { _3571,
                     _2082 };
    assign _2086 = _2083 + _2085;
    assign _2089 = _2086 + _2088;
    assign _2092 = _2089 + _2091;
    assign _2095 = _2092 + _2094;
    assign _2098 = _2095 + _2097;
    assign _2101 = _2098 + _2100;
    assign _2104 = _2101 + _2103;
    assign _2106 = _2104 < _3574;
    assign _2107 = _1770 & _2106;
    assign _3402 = ~ _2107;
    assign _3403 = _1770 & _3402;
    assign _3404 = _219 ? _3403 : _1770;
    assign _3405 = _529 ? _1800 : _3404;
    assign _159 = _3405;
    always @(posedge _207) begin
        if (_221)
            _1770 <= _2927;
        else
            _1770 <= _159;
    end
    assign _2124 = { _3571,
                     _1770 };
    assign _2121 = { _3571,
                     _1830 };
    assign _2118 = { _3571,
                     _2052 };
    assign _2115 = { _3571,
                     _2082 };
    assign _2113 = { _3571,
                     _2112 };
    assign _2116 = _2113 + _2115;
    assign _2119 = _2116 + _2118;
    assign _2122 = _2119 + _2121;
    assign _2125 = _2122 + _2124;
    assign _2128 = _2125 + _2127;
    assign _2131 = _2128 + _2130;
    assign _2134 = _2131 + _2133;
    assign _2136 = _2134 < _3574;
    assign _2137 = _1800 & _2136;
    assign _3406 = ~ _2137;
    assign _3407 = _1800 & _3406;
    assign _3408 = _219 ? _3407 : _1800;
    assign _3409 = _529 ? _1830 : _3408;
    assign _160 = _3409;
    always @(posedge _207) begin
        if (_221)
            _1800 <= _2927;
        else
            _1800 <= _160;
    end
    assign _2146 = { _3571,
                     _1800 };
    assign _2143 = { _3571,
                     _2082 };
    assign _2141 = { _3571,
                     _2112 };
    assign _2144 = _2141 + _2143;
    assign _2147 = _2144 + _2146;
    assign _2150 = _2147 + _2149;
    assign _2153 = _2150 + _2152;
    assign _2155 = _2153 < _3574;
    assign _2156 = _1830 & _2155;
    assign _3410 = ~ _2156;
    assign _3411 = _1830 & _3410;
    assign _3412 = _219 ? _3411 : _1830;
    assign _3413 = _529 ? _1883 : _3412;
    assign _161 = _3413;
    always @(posedge _207) begin
        if (_221)
            _1830 <= _2927;
        else
            _1830 <= _161;
    end
    assign _2431 = { _3571,
                     _1830 };
    assign _2428 = { _3571,
                     _2082 };
    assign _2425 = { _3571,
                     _2364 };
    assign _2423 = { _3571,
                     _2394 };
    assign _2426 = _2423 + _2425;
    assign _2429 = _2426 + _2428;
    assign _2432 = _2429 + _2431;
    assign _2435 = _2432 + _2434;
    assign _2437 = _2435 < _3574;
    assign _2438 = _2112 & _2437;
    assign _3414 = ~ _2438;
    assign _3415 = _2112 & _3414;
    assign _3416 = _219 ? _3415 : _2112;
    assign _3417 = _529 ? _2165 : _3416;
    assign _162 = _3417;
    always @(posedge _207) begin
        if (_221)
            _2112 <= _2927;
        else
            _2112 <= _162;
    end
    assign _2403 = { _3571,
                     _2112 };
    assign _2400 = { _3571,
                     _2334 };
    assign _2397 = { _3571,
                     _2364 };
    assign _2395 = { _3571,
                     _2394 };
    assign _2398 = _2395 + _2397;
    assign _2401 = _2398 + _2400;
    assign _2404 = _2401 + _2403;
    assign _2407 = _2404 + _2406;
    assign _2410 = _2407 + _2409;
    assign _2413 = _2410 + _2412;
    assign _2416 = _2413 + _2415;
    assign _2418 = _2416 < _3574;
    assign _2419 = _2082 & _2418;
    assign _3418 = ~ _2419;
    assign _3419 = _2082 & _3418;
    assign _3420 = _219 ? _3419 : _2082;
    assign _3421 = _529 ? _2112 : _3420;
    assign _163 = _3421;
    always @(posedge _207) begin
        if (_221)
            _2082 <= _2927;
        else
            _2082 <= _163;
    end
    assign _2373 = { _3571,
                     _2082 };
    assign _2370 = { _3571,
                     _2304 };
    assign _2367 = { _3571,
                     _2334 };
    assign _2365 = { _3571,
                     _2364 };
    assign _2368 = _2365 + _2367;
    assign _2371 = _2368 + _2370;
    assign _2374 = _2371 + _2373;
    assign _2377 = _2374 + _2376;
    assign _2380 = _2377 + _2379;
    assign _2383 = _2380 + _2382;
    assign _2386 = _2383 + _2385;
    assign _2388 = _2386 < _3574;
    assign _2389 = _2052 & _2388;
    assign _3422 = ~ _2389;
    assign _3423 = _2052 & _3422;
    assign _3424 = _219 ? _3423 : _2052;
    assign _3425 = _529 ? _2082 : _3424;
    assign _164 = _3425;
    always @(posedge _207) begin
        if (_221)
            _2052 <= _2927;
        else
            _2052 <= _164;
    end
    assign _2343 = { _3571,
                     _2052 };
    assign _2340 = { _3571,
                     _2274 };
    assign _2337 = { _3571,
                     _2304 };
    assign _2335 = { _3571,
                     _2334 };
    assign _2338 = _2335 + _2337;
    assign _2341 = _2338 + _2340;
    assign _2344 = _2341 + _2343;
    assign _2347 = _2344 + _2346;
    assign _2350 = _2347 + _2349;
    assign _2353 = _2350 + _2352;
    assign _2356 = _2353 + _2355;
    assign _2358 = _2356 < _3574;
    assign _2359 = _2022 & _2358;
    assign _3426 = ~ _2359;
    assign _3427 = _2022 & _3426;
    assign _3428 = _219 ? _3427 : _2022;
    assign _3429 = _529 ? _2052 : _3428;
    assign _165 = _3429;
    always @(posedge _207) begin
        if (_221)
            _2022 <= _2927;
        else
            _2022 <= _165;
    end
    assign _2313 = { _3571,
                     _2022 };
    assign _2310 = { _3571,
                     _2244 };
    assign _2307 = { _3571,
                     _2274 };
    assign _2305 = { _3571,
                     _2304 };
    assign _2308 = _2305 + _2307;
    assign _2311 = _2308 + _2310;
    assign _2314 = _2311 + _2313;
    assign _2317 = _2314 + _2316;
    assign _2320 = _2317 + _2319;
    assign _2323 = _2320 + _2322;
    assign _2326 = _2323 + _2325;
    assign _2328 = _2326 < _3574;
    assign _2329 = _1992 & _2328;
    assign _3430 = ~ _2329;
    assign _3431 = _1992 & _3430;
    assign _3432 = _219 ? _3431 : _1992;
    assign _3433 = _529 ? _2022 : _3432;
    assign _166 = _3433;
    always @(posedge _207) begin
        if (_221)
            _1992 <= _2927;
        else
            _1992 <= _166;
    end
    assign _2283 = { _3571,
                     _1992 };
    assign _2280 = { _3571,
                     _2214 };
    assign _2277 = { _3571,
                     _2244 };
    assign _2275 = { _3571,
                     _2274 };
    assign _2278 = _2275 + _2277;
    assign _2281 = _2278 + _2280;
    assign _2284 = _2281 + _2283;
    assign _2287 = _2284 + _2286;
    assign _2290 = _2287 + _2289;
    assign _2293 = _2290 + _2292;
    assign _2296 = _2293 + _2295;
    assign _2298 = _2296 < _3574;
    assign _2299 = _1962 & _2298;
    assign _3434 = ~ _2299;
    assign _3435 = _1962 & _3434;
    assign _3436 = _219 ? _3435 : _1962;
    assign _3437 = _529 ? _1992 : _3436;
    assign _167 = _3437;
    always @(posedge _207) begin
        if (_221)
            _1962 <= _2927;
        else
            _1962 <= _167;
    end
    assign _2253 = { _3571,
                     _1962 };
    assign _2250 = { _3571,
                     _2184 };
    assign _2247 = { _3571,
                     _2214 };
    assign _2245 = { _3571,
                     _2244 };
    assign _2248 = _2245 + _2247;
    assign _2251 = _2248 + _2250;
    assign _2254 = _2251 + _2253;
    assign _2257 = _2254 + _2256;
    assign _2260 = _2257 + _2259;
    assign _2263 = _2260 + _2262;
    assign _2266 = _2263 + _2265;
    assign _2268 = _2266 < _3574;
    assign _2269 = _1932 & _2268;
    assign _3438 = ~ _2269;
    assign _3439 = _1932 & _3438;
    assign _3440 = _219 ? _3439 : _1932;
    assign _3441 = _529 ? _1962 : _3440;
    assign _168 = _3441;
    always @(posedge _207) begin
        if (_221)
            _1932 <= _2927;
        else
            _1932 <= _168;
    end
    assign _2223 = { _3571,
                     _1932 };
    assign _2220 = { _3571,
                     _2161 };
    assign _2217 = { _3571,
                     _2184 };
    assign _2215 = { _3571,
                     _2214 };
    assign _2218 = _2215 + _2217;
    assign _2221 = _2218 + _2220;
    assign _2224 = _2221 + _2223;
    assign _2227 = _2224 + _2226;
    assign _2230 = _2227 + _2229;
    assign _2233 = _2230 + _2232;
    assign _2236 = _2233 + _2235;
    assign _2238 = _2236 < _3574;
    assign _2239 = _1902 & _2238;
    assign _3442 = ~ _2239;
    assign _3443 = _1902 & _3442;
    assign _3444 = _219 ? _3443 : _1902;
    assign _3445 = _529 ? _1932 : _3444;
    assign _169 = _3445;
    always @(posedge _207) begin
        if (_221)
            _1902 <= _2927;
        else
            _1902 <= _169;
    end
    assign _2193 = { _3571,
                     _1902 };
    assign _2190 = { _3571,
                     _2165 };
    assign _2187 = { _3571,
                     _2161 };
    assign _2185 = { _3571,
                     _2184 };
    assign _2188 = _2185 + _2187;
    assign _2191 = _2188 + _2190;
    assign _2194 = _2191 + _2193;
    assign _2197 = _2194 + _2196;
    assign _2200 = _2197 + _2199;
    assign _2203 = _2200 + _2202;
    assign _2206 = _2203 + _2205;
    assign _2208 = _2206 < _3574;
    assign _2209 = _1879 & _2208;
    assign _3446 = ~ _2209;
    assign _3447 = _1879 & _3446;
    assign _3448 = _219 ? _3447 : _1879;
    assign _3449 = _529 ? _1902 : _3448;
    assign _170 = _3449;
    always @(posedge _207) begin
        if (_221)
            _1879 <= _2927;
        else
            _1879 <= _170;
    end
    assign _2454 = { _3571,
                     _1879 };
    assign _2451 = { _3571,
                     _2161 };
    assign _2448 = { _3571,
                     _2447 };
    assign _2444 = { _3571,
                     _2443 };
    assign _2449 = _2444 + _2448;
    assign _2452 = _2449 + _2451;
    assign _2455 = _2452 + _2454;
    assign _2458 = _2455 + _2457;
    assign _2460 = _2458 < _3574;
    assign _2461 = _2165 & _2460;
    assign _3450 = ~ _2461;
    assign _3451 = _2165 & _3450;
    assign _3452 = _219 ? _3451 : _2165;
    assign _3453 = _529 ? _2161 : _3452;
    assign _171 = _3453;
    always @(posedge _207) begin
        if (_221)
            _2165 <= _2927;
        else
            _2165 <= _171;
    end
    assign _2739 = { _3571,
                     _2165 };
    assign _2736 = { _3571,
                     _2161 };
    assign _2733 = { _3571,
                     _2443 };
    assign _2730 = { _3571,
                     _2729 };
    assign _2726 = { _3571,
                     _2725 };
    assign _2731 = _2726 + _2730;
    assign _2734 = _2731 + _2733;
    assign _2737 = _2734 + _2736;
    assign _2740 = _2737 + _2739;
    assign _2742 = _2740 < _3574;
    assign _2743 = _2447 & _2742;
    assign _3454 = ~ _2743;
    assign _3455 = _2447 & _3454;
    assign _3456 = _219 ? _3455 : _2447;
    assign _3457 = _529 ? _2443 : _3456;
    assign _172 = _3457;
    always @(posedge _207) begin
        if (_221)
            _2447 <= _2927;
        else
            _2447 <= _172;
    end
    assign _2472 = { _3571,
                     _2447 };
    assign _2469 = { _3571,
                     _2443 };
    assign _2467 = { _3571,
                     _2466 };
    assign _2470 = _2467 + _2469;
    assign _2473 = _2470 + _2472;
    assign _2476 = _2473 + _2475;
    assign _2479 = _2476 + _2478;
    assign _2482 = _2479 + _2481;
    assign _2485 = _2482 + _2484;
    assign _2488 = _2485 + _2487;
    assign _2490 = _2488 < _3574;
    assign _2491 = _2161 & _2490;
    assign _3458 = ~ _2491;
    assign _3459 = _2161 & _3458;
    assign _3460 = _219 ? _3459 : _2161;
    assign _3461 = _529 ? _2184 : _3460;
    assign _173 = _3461;
    always @(posedge _207) begin
        if (_221)
            _2161 <= _2927;
        else
            _2161 <= _173;
    end
    assign _2508 = { _3571,
                     _2161 };
    assign _2505 = { _3571,
                     _2214 };
    assign _2502 = { _3571,
                     _2443 };
    assign _2499 = { _3571,
                     _2466 };
    assign _2497 = { _3571,
                     _2496 };
    assign _2500 = _2497 + _2499;
    assign _2503 = _2500 + _2502;
    assign _2506 = _2503 + _2505;
    assign _2509 = _2506 + _2508;
    assign _2512 = _2509 + _2511;
    assign _2515 = _2512 + _2514;
    assign _2518 = _2515 + _2517;
    assign _2520 = _2518 < _3574;
    assign _2521 = _2184 & _2520;
    assign _3462 = ~ _2521;
    assign _3463 = _2184 & _3462;
    assign _3464 = _219 ? _3463 : _2184;
    assign _3465 = _529 ? _2214 : _3464;
    assign _174 = _3465;
    always @(posedge _207) begin
        if (_221)
            _2184 <= _2927;
        else
            _2184 <= _174;
    end
    assign _2538 = { _3571,
                     _2184 };
    assign _2535 = { _3571,
                     _2244 };
    assign _2532 = { _3571,
                     _2466 };
    assign _2529 = { _3571,
                     _2496 };
    assign _2527 = { _3571,
                     _2526 };
    assign _2530 = _2527 + _2529;
    assign _2533 = _2530 + _2532;
    assign _2536 = _2533 + _2535;
    assign _2539 = _2536 + _2538;
    assign _2542 = _2539 + _2541;
    assign _2545 = _2542 + _2544;
    assign _2548 = _2545 + _2547;
    assign _2550 = _2548 < _3574;
    assign _2551 = _2214 & _2550;
    assign _3466 = ~ _2551;
    assign _3467 = _2214 & _3466;
    assign _3468 = _219 ? _3467 : _2214;
    assign _3469 = _529 ? _2244 : _3468;
    assign _175 = _3469;
    always @(posedge _207) begin
        if (_221)
            _2214 <= _2927;
        else
            _2214 <= _175;
    end
    assign _2568 = { _3571,
                     _2214 };
    assign _2565 = { _3571,
                     _2274 };
    assign _2562 = { _3571,
                     _2496 };
    assign _2559 = { _3571,
                     _2526 };
    assign _2557 = { _3571,
                     _2556 };
    assign _2560 = _2557 + _2559;
    assign _2563 = _2560 + _2562;
    assign _2566 = _2563 + _2565;
    assign _2569 = _2566 + _2568;
    assign _2572 = _2569 + _2571;
    assign _2575 = _2572 + _2574;
    assign _2578 = _2575 + _2577;
    assign _2580 = _2578 < _3574;
    assign _2581 = _2244 & _2580;
    assign _3470 = ~ _2581;
    assign _3471 = _2244 & _3470;
    assign _3472 = _219 ? _3471 : _2244;
    assign _3473 = _529 ? _2274 : _3472;
    assign _176 = _3473;
    always @(posedge _207) begin
        if (_221)
            _2244 <= _2927;
        else
            _2244 <= _176;
    end
    assign _2598 = { _3571,
                     _2244 };
    assign _2595 = { _3571,
                     _2304 };
    assign _2592 = { _3571,
                     _2526 };
    assign _2589 = { _3571,
                     _2556 };
    assign _2587 = { _3571,
                     _2586 };
    assign _2590 = _2587 + _2589;
    assign _2593 = _2590 + _2592;
    assign _2596 = _2593 + _2595;
    assign _2599 = _2596 + _2598;
    assign _2602 = _2599 + _2601;
    assign _2605 = _2602 + _2604;
    assign _2608 = _2605 + _2607;
    assign _2610 = _2608 < _3574;
    assign _2611 = _2274 & _2610;
    assign _3474 = ~ _2611;
    assign _3475 = _2274 & _3474;
    assign _3476 = _219 ? _3475 : _2274;
    assign _3477 = _529 ? _2304 : _3476;
    assign _177 = _3477;
    always @(posedge _207) begin
        if (_221)
            _2274 <= _2927;
        else
            _2274 <= _177;
    end
    assign _2628 = { _3571,
                     _2274 };
    assign _2625 = { _3571,
                     _2334 };
    assign _2622 = { _3571,
                     _2556 };
    assign _2619 = { _3571,
                     _2586 };
    assign _2617 = { _3571,
                     _2616 };
    assign _2620 = _2617 + _2619;
    assign _2623 = _2620 + _2622;
    assign _2626 = _2623 + _2625;
    assign _2629 = _2626 + _2628;
    assign _2632 = _2629 + _2631;
    assign _2635 = _2632 + _2634;
    assign _2638 = _2635 + _2637;
    assign _2640 = _2638 < _3574;
    assign _2641 = _2304 & _2640;
    assign _3478 = ~ _2641;
    assign _3479 = _2304 & _3478;
    assign _3480 = _219 ? _3479 : _2304;
    assign _3481 = _529 ? _2334 : _3480;
    assign _178 = _3481;
    always @(posedge _207) begin
        if (_221)
            _2304 <= _2927;
        else
            _2304 <= _178;
    end
    assign _2658 = { _3571,
                     _2304 };
    assign _2655 = { _3571,
                     _2364 };
    assign _2652 = { _3571,
                     _2586 };
    assign _2649 = { _3571,
                     _2616 };
    assign _2647 = { _3571,
                     _2646 };
    assign _2650 = _2647 + _2649;
    assign _2653 = _2650 + _2652;
    assign _2656 = _2653 + _2655;
    assign _2659 = _2656 + _2658;
    assign _2662 = _2659 + _2661;
    assign _2665 = _2662 + _2664;
    assign _2668 = _2665 + _2667;
    assign _2670 = _2668 < _3574;
    assign _2671 = _2334 & _2670;
    assign _3482 = ~ _2671;
    assign _3483 = _2334 & _3482;
    assign _3484 = _219 ? _3483 : _2334;
    assign _3485 = _529 ? _2364 : _3484;
    assign _179 = _3485;
    always @(posedge _207) begin
        if (_221)
            _2334 <= _2927;
        else
            _2334 <= _179;
    end
    assign _2688 = { _3571,
                     _2334 };
    assign _2685 = { _3571,
                     _2394 };
    assign _2682 = { _3571,
                     _2616 };
    assign _2679 = { _3571,
                     _2646 };
    assign _2677 = { _3571,
                     _2676 };
    assign _2680 = _2677 + _2679;
    assign _2683 = _2680 + _2682;
    assign _2686 = _2683 + _2685;
    assign _2689 = _2686 + _2688;
    assign _2692 = _2689 + _2691;
    assign _2695 = _2692 + _2694;
    assign _2698 = _2695 + _2697;
    assign _2700 = _2698 < _3574;
    assign _2701 = _2364 & _2700;
    assign _3486 = ~ _2701;
    assign _3487 = _2364 & _3486;
    assign _3488 = _219 ? _3487 : _2364;
    assign _3489 = _529 ? _2394 : _3488;
    assign _180 = _3489;
    always @(posedge _207) begin
        if (_221)
            _2364 <= _2927;
        else
            _2364 <= _180;
    end
    assign _2710 = { _3571,
                     _2364 };
    assign _2707 = { _3571,
                     _2646 };
    assign _2705 = { _3571,
                     _2676 };
    assign _2708 = _2705 + _2707;
    assign _2711 = _2708 + _2710;
    assign _2714 = _2711 + _2713;
    assign _2717 = _2714 + _2716;
    assign _2719 = _2717 < _3574;
    assign _2720 = _2394 & _2719;
    assign _3490 = ~ _2720;
    assign _3491 = _2394 & _3490;
    assign _3492 = _219 ? _3491 : _2394;
    assign _3493 = _529 ? _2447 : _3492;
    assign _181 = _3493;
    always @(posedge _207) begin
        if (_221)
            _2394 <= _2927;
        else
            _2394 <= _181;
    end
    assign _2995 = { _3571,
                     _2394 };
    assign _2992 = { _3571,
                     _2646 };
    assign _2989 = { _3571,
                     _2928 };
    assign _2987 = { _3571,
                     _2958 };
    assign _2990 = _2987 + _2989;
    assign _2993 = _2990 + _2992;
    assign _2996 = _2993 + _2995;
    assign _2999 = _2996 + _2998;
    assign _3001 = _2999 < _3574;
    assign _3002 = _2676 & _3001;
    assign _3494 = ~ _3002;
    assign _3495 = _2676 & _3494;
    assign _3496 = _219 ? _3495 : _2676;
    assign _3497 = _529 ? _2729 : _3496;
    assign _182 = _3497;
    always @(posedge _207) begin
        if (_221)
            _2676 <= _2927;
        else
            _2676 <= _182;
    end
    assign _2967 = { _3571,
                     _2676 };
    assign _2964 = { _3571,
                     _2898 };
    assign _2961 = { _3571,
                     _2928 };
    assign _2959 = { _3571,
                     _2958 };
    assign _2962 = _2959 + _2961;
    assign _2965 = _2962 + _2964;
    assign _2968 = _2965 + _2967;
    assign _2971 = _2968 + _2970;
    assign _2974 = _2971 + _2973;
    assign _2977 = _2974 + _2976;
    assign _2980 = _2977 + _2979;
    assign _2982 = _2980 < _3574;
    assign _2983 = _2646 & _2982;
    assign _3498 = ~ _2983;
    assign _3499 = _2646 & _3498;
    assign _3500 = _219 ? _3499 : _2646;
    assign _3501 = _529 ? _2676 : _3500;
    assign _183 = _3501;
    always @(posedge _207) begin
        if (_221)
            _2646 <= _2927;
        else
            _2646 <= _183;
    end
    assign _2937 = { _3571,
                     _2646 };
    assign _2934 = { _3571,
                     _2868 };
    assign _2931 = { _3571,
                     _2898 };
    assign _2929 = { _3571,
                     _2928 };
    assign _2932 = _2929 + _2931;
    assign _2935 = _2932 + _2934;
    assign _2938 = _2935 + _2937;
    assign _2941 = _2938 + _2940;
    assign _2944 = _2941 + _2943;
    assign _2947 = _2944 + _2946;
    assign _2950 = _2947 + _2949;
    assign _2952 = _2950 < _3574;
    assign _2953 = _2616 & _2952;
    assign _3502 = ~ _2953;
    assign _3503 = _2616 & _3502;
    assign _3504 = _219 ? _3503 : _2616;
    assign _3505 = _529 ? _2646 : _3504;
    assign _184 = _3505;
    always @(posedge _207) begin
        if (_221)
            _2616 <= _2927;
        else
            _2616 <= _184;
    end
    assign _2907 = { _3571,
                     _2616 };
    assign _2904 = { _3571,
                     _2838 };
    assign _2901 = { _3571,
                     _2868 };
    assign _2899 = { _3571,
                     _2898 };
    assign _2902 = _2899 + _2901;
    assign _2905 = _2902 + _2904;
    assign _2908 = _2905 + _2907;
    assign _2911 = _2908 + _2910;
    assign _2914 = _2911 + _2913;
    assign _2917 = _2914 + _2916;
    assign _2920 = _2917 + _2919;
    assign _2922 = _2920 < _3574;
    assign _2923 = _2586 & _2922;
    assign _3506 = ~ _2923;
    assign _3507 = _2586 & _3506;
    assign _3508 = _219 ? _3507 : _2586;
    assign _3509 = _529 ? _2616 : _3508;
    assign _185 = _3509;
    always @(posedge _207) begin
        if (_221)
            _2586 <= _2927;
        else
            _2586 <= _185;
    end
    assign _2877 = { _3571,
                     _2586 };
    assign _2874 = { _3571,
                     _2808 };
    assign _2871 = { _3571,
                     _2838 };
    assign _2869 = { _3571,
                     _2868 };
    assign _2872 = _2869 + _2871;
    assign _2875 = _2872 + _2874;
    assign _2878 = _2875 + _2877;
    assign _2881 = _2878 + _2880;
    assign _2884 = _2881 + _2883;
    assign _2887 = _2884 + _2886;
    assign _2890 = _2887 + _2889;
    assign _2892 = _2890 < _3574;
    assign _2893 = _2556 & _2892;
    assign _3510 = ~ _2893;
    assign _3511 = _2556 & _3510;
    assign _3512 = _219 ? _3511 : _2556;
    assign _3513 = _529 ? _2586 : _3512;
    assign _186 = _3513;
    always @(posedge _207) begin
        if (_221)
            _2556 <= _2927;
        else
            _2556 <= _186;
    end
    assign _2847 = { _3571,
                     _2556 };
    assign _2844 = { _3571,
                     _2778 };
    assign _2841 = { _3571,
                     _2808 };
    assign _2839 = { _3571,
                     _2838 };
    assign _2842 = _2839 + _2841;
    assign _2845 = _2842 + _2844;
    assign _2848 = _2845 + _2847;
    assign _2851 = _2848 + _2850;
    assign _2854 = _2851 + _2853;
    assign _2857 = _2854 + _2856;
    assign _2860 = _2857 + _2859;
    assign _2862 = _2860 < _3574;
    assign _2863 = _2526 & _2862;
    assign _3514 = ~ _2863;
    assign _3515 = _2526 & _3514;
    assign _3516 = _219 ? _3515 : _2526;
    assign _3517 = _529 ? _2556 : _3516;
    assign _187 = _3517;
    always @(posedge _207) begin
        if (_221)
            _2526 <= _2927;
        else
            _2526 <= _187;
    end
    assign _2817 = { _3571,
                     _2526 };
    assign _2814 = { _3571,
                     _2748 };
    assign _2811 = { _3571,
                     _2778 };
    assign _2809 = { _3571,
                     _2808 };
    assign _2812 = _2809 + _2811;
    assign _2815 = _2812 + _2814;
    assign _2818 = _2815 + _2817;
    assign _2821 = _2818 + _2820;
    assign _2824 = _2821 + _2823;
    assign _2827 = _2824 + _2826;
    assign _2830 = _2827 + _2829;
    assign _2832 = _2830 < _3574;
    assign _2833 = _2496 & _2832;
    assign _3518 = ~ _2833;
    assign _3519 = _2496 & _3518;
    assign _3520 = _219 ? _3519 : _2496;
    assign _3521 = _529 ? _2526 : _3520;
    assign _188 = _3521;
    always @(posedge _207) begin
        if (_221)
            _2496 <= _2927;
        else
            _2496 <= _188;
    end
    assign _2787 = { _3571,
                     _2496 };
    assign _2784 = { _3571,
                     _2725 };
    assign _2781 = { _3571,
                     _2748 };
    assign _2779 = { _3571,
                     _2778 };
    assign _2782 = _2779 + _2781;
    assign _2785 = _2782 + _2784;
    assign _2788 = _2785 + _2787;
    assign _2791 = _2788 + _2790;
    assign _2794 = _2791 + _2793;
    assign _2797 = _2794 + _2796;
    assign _2800 = _2797 + _2799;
    assign _2802 = _2800 < _3574;
    assign _2803 = _2466 & _2802;
    assign _3522 = ~ _2803;
    assign _3523 = _2466 & _3522;
    assign _3524 = _219 ? _3523 : _2466;
    assign _3525 = _529 ? _2496 : _3524;
    assign _189 = _3525;
    always @(posedge _207) begin
        if (_221)
            _2466 <= _2927;
        else
            _2466 <= _189;
    end
    assign _2757 = { _3571,
                     _2466 };
    assign _2754 = { _3571,
                     _2729 };
    assign _2751 = { _3571,
                     _2725 };
    assign _2749 = { _3571,
                     _2748 };
    assign _2752 = _2749 + _2751;
    assign _2755 = _2752 + _2754;
    assign _2758 = _2755 + _2757;
    assign _2761 = _2758 + _2760;
    assign _2764 = _2761 + _2763;
    assign _2767 = _2764 + _2766;
    assign _2770 = _2767 + _2769;
    assign _2772 = _2770 < _3574;
    assign _2773 = _2443 & _2772;
    assign _3526 = ~ _2773;
    assign _3527 = _2443 & _3526;
    assign _3528 = _219 ? _3527 : _2443;
    assign _3529 = _529 ? _2466 : _3528;
    assign _190 = _3529;
    always @(posedge _207) begin
        if (_221)
            _2443 <= _2927;
        else
            _2443 <= _190;
    end
    assign _3008 = { _3571,
                     _2443 };
    assign _3006 = { _3571,
                     _2725 };
    assign _3009 = _3006 + _3008;
    assign _3012 = _3009 + _3011;
    assign _3014 = _3012 < _3574;
    assign _3015 = _2729 & _3014;
    assign _3530 = ~ _3015;
    assign _3531 = _2729 & _3530;
    assign _3532 = _219 ? _3531 : _2729;
    assign _3533 = _529 ? _2725 : _3532;
    assign _191 = _3533;
    always @(posedge _207) begin
        if (_221)
            _2729 <= _2927;
        else
            _2729 <= _191;
    end
    assign _3021 = { _3571,
                     _2729 };
    assign _3019 = { _3571,
                     _2748 };
    assign _3022 = _3019 + _3021;
    assign _3025 = _3022 + _3024;
    assign _3028 = _3025 + _3027;
    assign _3031 = _3028 + _3030;
    assign _3033 = _3031 < _3574;
    assign _3034 = _2725 & _3033;
    assign _3534 = ~ _3034;
    assign _3535 = _2725 & _3534;
    assign _3536 = _219 ? _3535 : _2725;
    assign _3537 = _529 ? _2748 : _3536;
    assign _192 = _3537;
    always @(posedge _207) begin
        if (_221)
            _2725 <= _2927;
        else
            _2725 <= _192;
    end
    assign _3040 = { _3571,
                     _2725 };
    assign _3038 = { _3571,
                     _2778 };
    assign _3041 = _3038 + _3040;
    assign _3044 = _3041 + _3043;
    assign _3047 = _3044 + _3046;
    assign _3050 = _3047 + _3049;
    assign _3052 = _3050 < _3574;
    assign _3053 = _2748 & _3052;
    assign _3538 = ~ _3053;
    assign _3539 = _2748 & _3538;
    assign _3540 = _219 ? _3539 : _2748;
    assign _3541 = _529 ? _2778 : _3540;
    assign _193 = _3541;
    always @(posedge _207) begin
        if (_221)
            _2748 <= _2927;
        else
            _2748 <= _193;
    end
    assign _3059 = { _3571,
                     _2748 };
    assign _3057 = { _3571,
                     _2808 };
    assign _3060 = _3057 + _3059;
    assign _3063 = _3060 + _3062;
    assign _3066 = _3063 + _3065;
    assign _3069 = _3066 + _3068;
    assign _3071 = _3069 < _3574;
    assign _3072 = _2778 & _3071;
    assign _3542 = ~ _3072;
    assign _3543 = _2778 & _3542;
    assign _3544 = _219 ? _3543 : _2778;
    assign _3545 = _529 ? _2808 : _3544;
    assign _194 = _3545;
    always @(posedge _207) begin
        if (_221)
            _2778 <= _2927;
        else
            _2778 <= _194;
    end
    assign _3078 = { _3571,
                     _2778 };
    assign _3076 = { _3571,
                     _2838 };
    assign _3079 = _3076 + _3078;
    assign _3082 = _3079 + _3081;
    assign _3085 = _3082 + _3084;
    assign _3088 = _3085 + _3087;
    assign _3090 = _3088 < _3574;
    assign _3091 = _2808 & _3090;
    assign _3546 = ~ _3091;
    assign _3547 = _2808 & _3546;
    assign _3548 = _219 ? _3547 : _2808;
    assign _3549 = _529 ? _2838 : _3548;
    assign _195 = _3549;
    always @(posedge _207) begin
        if (_221)
            _2808 <= _2927;
        else
            _2808 <= _195;
    end
    assign _3097 = { _3571,
                     _2808 };
    assign _3095 = { _3571,
                     _2868 };
    assign _3098 = _3095 + _3097;
    assign _3101 = _3098 + _3100;
    assign _3104 = _3101 + _3103;
    assign _3107 = _3104 + _3106;
    assign _3109 = _3107 < _3574;
    assign _3110 = _2838 & _3109;
    assign _3550 = ~ _3110;
    assign _3551 = _2838 & _3550;
    assign _3552 = _219 ? _3551 : _2838;
    assign _3553 = _529 ? _2868 : _3552;
    assign _196 = _3553;
    always @(posedge _207) begin
        if (_221)
            _2838 <= _2927;
        else
            _2838 <= _196;
    end
    assign _3116 = { _3571,
                     _2838 };
    assign _3114 = { _3571,
                     _2898 };
    assign _3117 = _3114 + _3116;
    assign _3120 = _3117 + _3119;
    assign _3123 = _3120 + _3122;
    assign _3126 = _3123 + _3125;
    assign _3128 = _3126 < _3574;
    assign _3129 = _2868 & _3128;
    assign _3554 = ~ _3129;
    assign _3555 = _2868 & _3554;
    assign _3556 = _219 ? _3555 : _2868;
    assign _3557 = _529 ? _2898 : _3556;
    assign _197 = _3557;
    always @(posedge _207) begin
        if (_221)
            _2868 <= _2927;
        else
            _2868 <= _197;
    end
    assign _3135 = { _3571,
                     _2868 };
    assign _3133 = { _3571,
                     _2928 };
    assign _3136 = _3133 + _3135;
    assign _3139 = _3136 + _3138;
    assign _3142 = _3139 + _3141;
    assign _3145 = _3142 + _3144;
    assign _3147 = _3145 < _3574;
    assign _3148 = _2898 & _3147;
    assign _3558 = ~ _3148;
    assign _3559 = _2898 & _3558;
    assign _3560 = _219 ? _3559 : _2898;
    assign _3561 = _529 ? _2928 : _3560;
    assign _198 = _3561;
    always @(posedge _207) begin
        if (_221)
            _2898 <= _2927;
        else
            _2898 <= _198;
    end
    assign _3154 = { _3571,
                     _2898 };
    assign _3152 = { _3571,
                     _2958 };
    assign _3155 = _3152 + _3154;
    assign _3158 = _3155 + _3157;
    assign _3161 = _3158 + _3160;
    assign _3164 = _3161 + _3163;
    assign _3166 = _3164 < _3574;
    assign _3167 = _2928 & _3166;
    assign _3562 = ~ _3167;
    assign _3563 = _2928 & _3562;
    assign _3564 = _219 ? _3563 : _2928;
    assign _3565 = _529 ? _2958 : _3564;
    assign _199 = _3565;
    always @(posedge _207) begin
        if (_221)
            _2928 <= _2927;
        else
            _2928 <= _199;
    end
    assign _3567 = { _3571,
                     _2928 };
    assign _3570 = _3567 + _3569;
    assign _3573 = _3570 + _3572;
    assign _3575 = _3573 < _3574;
    assign _220 = _218[1:1];
    assign _221 = _205 | _220;
    assign _3580 = _209[0:0];
    assign _3577 = ~ _3576;
    assign _3578 = _2958 & _3577;
    assign _3579 = _219 ? _3578 : _2958;
    assign _3581 = _529 ? _3580 : _3579;
    assign _200 = _3581;
    always @(posedge _207) begin
        if (_221)
            _2958 <= _2927;
        else
            _2958 <= _200;
    end
    assign _3576 = _2958 & _3575;
    assign gnd = 1'b0;
    assign _3582 = _219 ? _3576 : gnd;
    assign _527 = 4'b0001;
    assign _528 = _212 == _527;
    assign _529 = _203 & _528;
    assign _3583 = _529 ? gnd : _3582;
    assign _201 = _3583;
    assign _227 = { _3889,
                    _201 };
    assign _230 = _227 + _229;
    assign _233 = _230 + _232;
    assign _236 = _233 + _235;
    assign _239 = _236 + _238;
    assign _242 = _239 + _241;
    assign _245 = _242 + _244;
    assign _248 = _245 + _247;
    assign _251 = _248 + _250;
    assign _254 = _251 + _253;
    assign _257 = _254 + _256;
    assign _260 = _257 + _259;
    assign _263 = _260 + _262;
    assign _266 = _263 + _265;
    assign _269 = _266 + _268;
    assign _272 = _269 + _271;
    assign _275 = _272 + _274;
    assign _278 = _275 + _277;
    assign _281 = _278 + _280;
    assign _284 = _281 + _283;
    assign _287 = _284 + _286;
    assign _290 = _287 + _289;
    assign _293 = _290 + _292;
    assign _296 = _293 + _295;
    assign _299 = _296 + _298;
    assign _302 = _299 + _301;
    assign _305 = _302 + _304;
    assign _308 = _305 + _307;
    assign _311 = _308 + _310;
    assign _314 = _311 + _313;
    assign _317 = _314 + _316;
    assign _320 = _317 + _319;
    assign _323 = _320 + _322;
    assign _326 = _323 + _325;
    assign _329 = _326 + _328;
    assign _332 = _329 + _331;
    assign _335 = _332 + _334;
    assign _338 = _335 + _337;
    assign _341 = _338 + _340;
    assign _344 = _341 + _343;
    assign _347 = _344 + _346;
    assign _350 = _347 + _349;
    assign _353 = _350 + _352;
    assign _356 = _353 + _355;
    assign _359 = _356 + _358;
    assign _362 = _359 + _361;
    assign _365 = _362 + _364;
    assign _368 = _365 + _367;
    assign _371 = _368 + _370;
    assign _374 = _371 + _373;
    assign _377 = _374 + _376;
    assign _380 = _377 + _379;
    assign _383 = _380 + _382;
    assign _386 = _383 + _385;
    assign _389 = _386 + _388;
    assign _392 = _389 + _391;
    assign _395 = _392 + _394;
    assign _398 = _395 + _397;
    assign _401 = _398 + _400;
    assign _404 = _401 + _403;
    assign _407 = _404 + _406;
    assign _410 = _407 + _409;
    assign _413 = _410 + _412;
    assign _416 = _413 + _415;
    assign _419 = _416 + _418;
    assign _422 = _419 + _421;
    assign _425 = _422 + _424;
    assign _428 = _425 + _427;
    assign _431 = _428 + _430;
    assign _434 = _431 + _433;
    assign _437 = _434 + _436;
    assign _440 = _437 + _439;
    assign _443 = _440 + _442;
    assign _446 = _443 + _445;
    assign _449 = _446 + _448;
    assign _452 = _449 + _451;
    assign _455 = _452 + _454;
    assign _458 = _455 + _457;
    assign _461 = _458 + _460;
    assign _464 = _461 + _463;
    assign _467 = _464 + _466;
    assign _470 = _467 + _469;
    assign _473 = _470 + _472;
    assign _476 = _473 + _475;
    assign _479 = _476 + _478;
    assign _482 = _479 + _481;
    assign _485 = _482 + _484;
    assign _488 = _485 + _487;
    assign _491 = _488 + _490;
    assign _494 = _491 + _493;
    assign _497 = _494 + _496;
    assign _500 = _497 + _499;
    assign _503 = _500 + _502;
    assign _506 = _503 + _505;
    assign _509 = _506 + _508;
    assign _512 = _509 + _511;
    assign _515 = _512 + _514;
    assign _518 = _515 + _517;
    assign _521 = _518 + _520;
    assign _524 = _521 + _523;
    assign _3587 = _524 == _3592;
    assign _219 = _218[0:0];
    assign _3588 = _219 & _3587;
    assign _3585 = 31'b0000000000000000000000000000000;
    assign _3589 = { _3585,
                     _3588 };
    assign _3584 = 32'b00000000000000000000000000000000;
    assign _215 = 4'b0000;
    assign _216 = _212 == _215;
    assign _203 = write_enable;
    assign _217 = _203 & _216;
    assign _205 = clear;
    assign _207 = clock;
    assign _209 = write_data;
    assign _210 = _209;
    always @(posedge _207) begin
        if (_205)
            _218 <= _3584;
        else
            if (_217)
                _218 <= _210;
    end
    assign _212 = write_addr;
    always @* begin
        case (_212)
        0:
            _3893 <= _218;
        1:
            _3893 <= _3584;
        2:
            _3893 <= _3589;
        3:
            _3893 <= _3591;
        default:
            _3893 <= _3892;
        endcase
    end
    assign read_data = _3893;

endmodule
module aoc_solver_top (
    write_data,
    write_addr,
    write_enable,
    clear,
    clock,
    read_data
);

    input [31:0] write_data;
    input [3:0] write_addr;
    input write_enable;
    input clear;
    input clock;
    output [31:0] read_data;

    wire [31:0] _2;
    wire [3:0] _4;
    wire _6;
    wire _8;
    wire _10;
    wire [31:0] _13;
    wire [31:0] _11;
    assign _2 = write_data;
    assign _4 = write_addr;
    assign _6 = write_enable;
    assign _8 = clear;
    assign _10 = clock;
    aoc_solver
        aoc_solver
        ( .clock(_10),
          .clear(_8),
          .write_enable(_6),
          .write_addr(_4),
          .write_data(_2),
          .read_data(_13[31:0]) );
    assign _11 = _13;
    assign read_data = _11;

endmodule

